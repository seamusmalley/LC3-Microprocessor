<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-152.367,32.0587,315.996,-209.762</PageViewport>
<gate>
<ID>389</ID>
<type>EE_VDD</type>
<position>2,-117.5</position>
<output>
<ID>OUT_0</ID>395 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>391</ID>
<type>EE_VDD</type>
<position>9.5,-117.5</position>
<output>
<ID>OUT_0</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_REGISTER8</type>
<position>0.5,-165</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>84 </input>
<output>
<ID>OUT_0</ID>11 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>30 </output>
<output>
<ID>OUT_4</ID>29 </output>
<output>
<ID>OUT_5</ID>28 </output>
<output>
<ID>OUT_6</ID>27 </output>
<output>
<ID>OUT_7</ID>26 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>385 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>-112.5,50</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>-112.5,43.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>-80.5,-155</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-80,-148.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>15.5,-163.5</position>
<gparam>LABEL_TEXT LD.MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>1,-158.5</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AE_REGISTER8</type>
<position>-37.5,-165</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>47 </input>
<input>
<ID>IN_3</ID>48 </input>
<input>
<ID>IN_4</ID>49 </input>
<input>
<ID>IN_5</ID>50 </input>
<input>
<ID>IN_6</ID>51 </input>
<input>
<ID>IN_7</ID>52 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>41 </output>
<output>
<ID>OUT_2</ID>42 </output>
<output>
<ID>OUT_3</ID>43 </output>
<output>
<ID>OUT_4</ID>44 </output>
<output>
<ID>OUT_5</ID>36 </output>
<output>
<ID>OUT_6</ID>37 </output>
<output>
<ID>OUT_7</ID>38 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>5 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-53,-165.5</position>
<gparam>LABEL_TEXT LD.MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>1,-197</position>
<gparam>LABEL_TEXT MEM.EN R,W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>15,-184</position>
<gparam>LABEL_TEXT MEMORY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-38,-159</position>
<input>
<ID>ENABLE_0</ID>53 </input>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>43 </input>
<input>
<ID>IN_4</ID>44 </input>
<input>
<ID>IN_5</ID>36 </input>
<input>
<ID>IN_6</ID>37 </input>
<input>
<ID>IN_7</ID>38 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>98 </output>
<output>
<ID>OUT_2</ID>97 </output>
<output>
<ID>OUT_3</ID>96 </output>
<output>
<ID>OUT_4</ID>95 </output>
<output>
<ID>OUT_5</ID>94 </output>
<output>
<ID>OUT_6</ID>93 </output>
<output>
<ID>OUT_7</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>-54,-159</position>
<gparam>LABEL_TEXT GateMDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>HA_JUNC_2</type>
<position>-107.5,49.5</position>
<input>
<ID>N_in1</ID>84 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>-47,-144.5</position>
<gparam>LABEL_TEXT LD.IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-156</position>
<input>
<ID>N_in1</ID>84 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>-14,-128</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>9,-127.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>33</ID>
<type>HA_JUNC_2</type>
<position>-107.5,48.5</position>
<input>
<ID>N_in1</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-155</position>
<input>
<ID>N_in1</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>HA_JUNC_2</type>
<position>-107.5,47.5</position>
<input>
<ID>N_in1</ID>94 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-154</position>
<input>
<ID>N_in1</ID>94 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>HA_JUNC_2</type>
<position>-107.5,46.5</position>
<input>
<ID>N_in1</ID>95 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-153</position>
<input>
<ID>N_in1</ID>95 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>HA_JUNC_2</type>
<position>-107.5,45.5</position>
<input>
<ID>N_in1</ID>96 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-152</position>
<input>
<ID>N_in1</ID>96 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>HA_JUNC_2</type>
<position>-107.5,44.5</position>
<input>
<ID>N_in1</ID>97 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-151</position>
<input>
<ID>N_in1</ID>97 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>HA_JUNC_2</type>
<position>-107.5,43.5</position>
<input>
<ID>N_in1</ID>98 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-150</position>
<input>
<ID>N_in1</ID>98 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>HA_JUNC_2</type>
<position>-107.5,42.5</position>
<input>
<ID>N_in1</ID>99 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>HA_JUNC_2</type>
<position>-74.5,-149</position>
<input>
<ID>N_in1</ID>99 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>8,-70.5</position>
<gparam>LABEL_TEXT BEN</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>52</ID>
<type>AE_RAM_8x8</type>
<position>0.5,-185</position>
<input>
<ID>ADDRESS_0</ID>11 </input>
<input>
<ID>ADDRESS_1</ID>32 </input>
<input>
<ID>ADDRESS_2</ID>31 </input>
<input>
<ID>ADDRESS_3</ID>30 </input>
<input>
<ID>ADDRESS_4</ID>29 </input>
<input>
<ID>ADDRESS_5</ID>28 </input>
<input>
<ID>ADDRESS_6</ID>27 </input>
<input>
<ID>ADDRESS_7</ID>26 </input>
<input>
<ID>DATA_IN_0</ID>9 </input>
<input>
<ID>DATA_IN_1</ID>8 </input>
<input>
<ID>DATA_IN_2</ID>7 </input>
<input>
<ID>DATA_IN_3</ID>6 </input>
<input>
<ID>DATA_IN_4</ID>4 </input>
<input>
<ID>DATA_IN_5</ID>3 </input>
<input>
<ID>DATA_IN_6</ID>2 </input>
<input>
<ID>DATA_IN_7</ID>1 </input>
<output>
<ID>DATA_OUT_0</ID>9 </output>
<output>
<ID>DATA_OUT_1</ID>8 </output>
<output>
<ID>DATA_OUT_2</ID>7 </output>
<output>
<ID>DATA_OUT_3</ID>6 </output>
<output>
<ID>DATA_OUT_4</ID>4 </output>
<output>
<ID>DATA_OUT_5</ID>3 </output>
<output>
<ID>DATA_OUT_6</ID>2 </output>
<output>
<ID>DATA_OUT_7</ID>1 </output>
<input>
<ID>ENABLE_0</ID>57 </input>
<input>
<ID>write_clock</ID>12 </input>
<input>
<ID>write_enable</ID>54 </input>
<gparam>angle 270</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>56</ID>
<type>AE_REGISTER8</type>
<position>-30,-144</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>84 </input>
<output>
<ID>OUT_0</ID>120 </output>
<output>
<ID>OUT_1</ID>121 </output>
<output>
<ID>OUT_2</ID>122 </output>
<output>
<ID>OUT_3</ID>119 </output>
<output>
<ID>OUT_4</ID>118 </output>
<output>
<ID>OUT_5</ID>117 </output>
<output>
<ID>OUT_6</ID>81 </output>
<output>
<ID>OUT_7</ID>80 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>21 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_REGISTER8</type>
<position>-18,-21</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<input>
<ID>IN_2</ID>209 </input>
<input>
<ID>IN_3</ID>210 </input>
<input>
<ID>IN_4</ID>211 </input>
<input>
<ID>IN_5</ID>212 </input>
<input>
<ID>IN_6</ID>213 </input>
<input>
<ID>IN_7</ID>214 </input>
<output>
<ID>OUT_0</ID>16 </output>
<output>
<ID>OUT_1</ID>17 </output>
<output>
<ID>OUT_2</ID>18 </output>
<output>
<ID>OUT_3</ID>19 </output>
<output>
<ID>OUT_4</ID>20 </output>
<output>
<ID>OUT_5</ID>13 </output>
<output>
<ID>OUT_6</ID>14 </output>
<output>
<ID>OUT_7</ID>15 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>22 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>62</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-18.5,-12</position>
<input>
<ID>ENABLE_0</ID>23 </input>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>19 </input>
<input>
<ID>IN_4</ID>20 </input>
<input>
<ID>IN_5</ID>13 </input>
<input>
<ID>IN_6</ID>14 </input>
<input>
<ID>IN_7</ID>15 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>98 </output>
<output>
<ID>OUT_2</ID>97 </output>
<output>
<ID>OUT_3</ID>96 </output>
<output>
<ID>OUT_4</ID>95 </output>
<output>
<ID>OUT_5</ID>94 </output>
<output>
<ID>OUT_6</ID>93 </output>
<output>
<ID>OUT_7</ID>84 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>31,-89.5</position>
<gparam>LABEL_TEXT COND + IRD</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>73</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-16,-185.5</position>
<input>
<ID>ENABLE_0</ID>54 </input>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>84 </input>
<output>
<ID>OUT_0</ID>9 </output>
<output>
<ID>OUT_1</ID>8 </output>
<output>
<ID>OUT_2</ID>7 </output>
<output>
<ID>OUT_3</ID>6 </output>
<output>
<ID>OUT_4</ID>4 </output>
<output>
<ID>OUT_5</ID>3 </output>
<output>
<ID>OUT_6</ID>2 </output>
<output>
<ID>OUT_7</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_MUX_2x1</type>
<position>-7,-120.5</position>
<input>
<ID>IN_0</ID>382 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>60 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_OR2</type>
<position>2,-111.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_MUX_2x1</type>
<position>1,-120.5</position>
<input>
<ID>IN_0</ID>394 </input>
<input>
<ID>IN_1</ID>395 </input>
<output>
<ID>OUT</ID>61 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_MUX_2x1</type>
<position>8.5,-120.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>396 </input>
<output>
<ID>OUT</ID>66 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_MUX_2x1</type>
<position>-13.5,-120.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>59 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_AND8</type>
<position>-49,-115</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<input>
<ID>IN_2</ID>88 </input>
<input>
<ID>IN_3</ID>87 </input>
<input>
<ID>IN_4</ID>89 </input>
<input>
<ID>IN_5</ID>90 </input>
<input>
<ID>IN_6</ID>91 </input>
<input>
<ID>IN_7</ID>92 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_OR2</type>
<position>-12.5,-112</position>
<input>
<ID>IN_0</ID>376 </input>
<input>
<ID>IN_1</ID>375 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>-51,-106</position>
<input>
<ID>N_in0</ID>84 </input>
<input>
<ID>N_in1</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-51,-103</position>
<gparam>LABEL_TEXT n</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-111.5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-112.5</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-113.5</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-114.5</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-115.5</position>
<input>
<ID>IN_0</ID>96 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-116.5</position>
<input>
<ID>IN_0</ID>97 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-117.5</position>
<input>
<ID>IN_0</ID>98 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_SMALL_INVERTER</type>
<position>-54,-118.5</position>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>95</ID>
<type>GA_LED</type>
<position>-45,-115</position>
<input>
<ID>N_in0</ID>100 </input>
<input>
<ID>N_in1</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>-45,-112</position>
<gparam>LABEL_TEXT z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND2</type>
<position>-30,-110.5</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_SMALL_INVERTER</type>
<position>-35,-109.5</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_SMALL_INVERTER</type>
<position>-35,-111.5</position>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>-22,-105</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>-26,-106.5</position>
<gparam>LABEL_TEXT p</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AF_DFF_LOW</type>
<position>-54.5,-81</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>110 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>clock_enable</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>-56.5,-75</position>
<gparam>LABEL_TEXT n</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>-41,-74.5</position>
<gparam>LABEL_TEXT z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>-28,-74.5</position>
<gparam>LABEL_TEXT p</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>-70.5,-78.5</position>
<gparam>LABEL_TEXT LD.CC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>GA_LED</type>
<position>-53,-75.5</position>
<input>
<ID>N_in1</ID>110 </input>
<input>
<ID>N_in3</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>-39,-75.5</position>
<input>
<ID>N_in1</ID>107 </input>
<input>
<ID>N_in3</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>GA_LED</type>
<position>-25.5,-75.5</position>
<input>
<ID>N_in1</ID>106 </input>
<input>
<ID>N_in3</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AF_DFF_LOW</type>
<position>-39.5,-81</position>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>107 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>clock_enable</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>114</ID>
<type>AF_DFF_LOW</type>
<position>-26,-81</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>106 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>clock_enable</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>-53,-65.5</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>-39.5,-65.5</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_AND2</type>
<position>-26,-65.5</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR3</type>
<position>2.5,-75.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<input>
<ID>IN_2</ID>116 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_REGISTER4</type>
<position>30,-79.5</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>137 </input>
<input>
<ID>IN_2</ID>138 </input>
<input>
<ID>IN_3</ID>139 </input>
<output>
<ID>OUT_0</ID>78 </output>
<output>
<ID>OUT_1</ID>63 </output>
<output>
<ID>OUT_2</ID>382 </output>
<output>
<ID>OUT_3</ID>376 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>142 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>123</ID>
<type>EE_VDD</type>
<position>36,-78.5</position>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_REGISTER4</type>
<position>30,-98.5</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_2</ID>145 </input>
<input>
<ID>IN_3</ID>147 </input>
<output>
<ID>OUT_0</ID>40 </output>
<output>
<ID>OUT_1</ID>79 </output>
<output>
<ID>OUT_2</ID>411 </output>
<output>
<ID>OUT_3</ID>377 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>179 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>125</ID>
<type>BA_ROM_4x4</type>
<position>30,-128</position>
<input>
<ID>ADDRESS_0</ID>66 </input>
<input>
<ID>ADDRESS_1</ID>61 </input>
<input>
<ID>ADDRESS_2</ID>60 </input>
<input>
<ID>ADDRESS_3</ID>59 </input>
<output>
<ID>DATA_OUT_0</ID>187 </output>
<output>
<ID>DATA_OUT_1</ID>196 </output>
<output>
<ID>DATA_OUT_2</ID>198 </output>
<output>
<ID>DATA_OUT_3</ID>188 </output>
<input>
<ID>ENABLE_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 8</lparam>
<lparam>Address:2 8</lparam>
<lparam>Address:8 6</lparam>
<lparam>Address:11 6</lparam>
<lparam>Address:12 1</lparam>
<lparam>Address:15 6</lparam></gate>
<gate>
<ID>127</ID>
<type>BA_ROM_4x4</type>
<position>30.5,-69</position>
<input>
<ID>ADDRESS_0</ID>66 </input>
<input>
<ID>ADDRESS_1</ID>61 </input>
<input>
<ID>ADDRESS_2</ID>60 </input>
<input>
<ID>ADDRESS_3</ID>59 </input>
<output>
<ID>DATA_OUT_0</ID>136 </output>
<output>
<ID>DATA_OUT_1</ID>137 </output>
<output>
<ID>DATA_OUT_2</ID>138 </output>
<output>
<ID>DATA_OUT_3</ID>139 </output>
<input>
<ID>ENABLE_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 10</lparam>
<lparam>Address:1 5</lparam>
<lparam>Address:3 4</lparam>
<lparam>Address:5 8</lparam>
<lparam>Address:7 1</lparam>
<lparam>Address:9 14</lparam>
<lparam>Address:10 12</lparam>
<lparam>Address:12 13</lparam>
<lparam>Address:14 6</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>-76,-57</position>
<gparam>LABEL_TEXT SEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>BA_ROM_4x4</type>
<position>30.5,-88.5</position>
<input>
<ID>ADDRESS_0</ID>66 </input>
<input>
<ID>ADDRESS_1</ID>61 </input>
<input>
<ID>ADDRESS_2</ID>60 </input>
<input>
<ID>ADDRESS_3</ID>59 </input>
<output>
<ID>DATA_OUT_0</ID>143 </output>
<output>
<ID>DATA_OUT_1</ID>144 </output>
<output>
<ID>DATA_OUT_2</ID>145 </output>
<output>
<ID>DATA_OUT_3</ID>147 </output>
<input>
<ID>ENABLE_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:4 2</lparam>
<lparam>Address:7 8</lparam>
<lparam>Address:13 1</lparam>
<lparam>Address:14 4</lparam></gate>
<gate>
<ID>130</ID>
<type>EE_VDD</type>
<position>36,-97.5</position>
<output>
<ID>OUT_0</ID>179 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>131</ID>
<type>BA_ROM_4x4</type>
<position>30,-108.5</position>
<input>
<ID>ADDRESS_0</ID>66 </input>
<input>
<ID>ADDRESS_1</ID>61 </input>
<input>
<ID>ADDRESS_2</ID>60 </input>
<input>
<ID>ADDRESS_3</ID>59 </input>
<output>
<ID>DATA_OUT_0</ID>182 </output>
<output>
<ID>DATA_OUT_1</ID>183 </output>
<output>
<ID>DATA_OUT_2</ID>184 </output>
<output>
<ID>DATA_OUT_3</ID>181 </output>
<input>
<ID>ENABLE_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 4</lparam>
<lparam>Address:1 8</lparam>
<lparam>Address:8 1</lparam>
<lparam>Address:9 8</lparam>
<lparam>Address:11 2</lparam>
<lparam>Address:12 1</lparam>
<lparam>Address:15 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_REGISTER4</type>
<position>29.5,-118</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>183 </input>
<input>
<ID>IN_2</ID>184 </input>
<input>
<ID>IN_3</ID>181 </input>
<output>
<ID>OUT_0</ID>53 </output>
<output>
<ID>OUT_1</ID>373 </output>
<output>
<ID>OUT_2</ID>23 </output>
<output>
<ID>OUT_3</ID>217 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>180 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>29,-77</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>134</ID>
<type>EE_VDD</type>
<position>35.5,-117</position>
<output>
<ID>OUT_0</ID>180 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_REGISTER4</type>
<position>30,-138</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>196 </input>
<input>
<ID>IN_2</ID>198 </input>
<input>
<ID>IN_3</ID>188 </input>
<output>
<ID>OUT_0</ID>21 </output>
<output>
<ID>OUT_1</ID>109 </output>
<output>
<ID>OUT_2</ID>264 </output>
<output>
<ID>OUT_3</ID>22 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>215 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>136</ID>
<type>EE_VDD</type>
<position>36,-137</position>
<output>
<ID>OUT_0</ID>215 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_AND2</type>
<position>3,-105.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_REGISTER4</type>
<position>54,-98</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>221 </input>
<input>
<ID>IN_3</ID>218 </input>
<output>
<ID>OUT_0</ID>54 </output>
<output>
<ID>OUT_1</ID>57 </output>
<output>
<ID>OUT_2</ID>5 </output>
<output>
<ID>OUT_3</ID>385 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>222 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>139</ID>
<type>EE_VDD</type>
<position>60,-97</position>
<output>
<ID>OUT_0</ID>222 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_REGISTER4</type>
<position>54,-120</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>322 </input>
<input>
<ID>IN_2</ID>383 </input>
<input>
<ID>IN_3</ID>269 </input>
<output>
<ID>OUT_0</ID>419 </output>
<output>
<ID>OUT_1</ID>185 </output>
<output>
<ID>OUT_2</ID>372 </output>
<output>
<ID>OUT_3</ID>141 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>384 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>141</ID>
<type>EE_VDD</type>
<position>60,-117.5</position>
<output>
<ID>OUT_0</ID>384 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>-81,-55</position>
<input>
<ID>N_in2</ID>122 </input>
<input>
<ID>N_in3</ID>160 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>GA_LED</type>
<position>-77.5,-55</position>
<input>
<ID>N_in2</ID>122 </input>
<input>
<ID>N_in3</ID>159 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>GA_LED</type>
<position>-74,-55</position>
<input>
<ID>N_in2</ID>122 </input>
<input>
<ID>N_in3</ID>158 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>GA_LED</type>
<position>-71,-55</position>
<input>
<ID>N_in2</ID>122 </input>
<input>
<ID>N_in3</ID>157 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>-68,-55</position>
<input>
<ID>N_in2</ID>122 </input>
<input>
<ID>N_in3</ID>156 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>-65,-55</position>
<input>
<ID>N_in2</ID>122 </input>
<input>
<ID>N_in3</ID>155 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>-62,-55</position>
<input>
<ID>N_in2</ID>121 </input>
<input>
<ID>N_in3</ID>154 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>-59,-55</position>
<input>
<ID>N_in2</ID>120 </input>
<input>
<ID>N_in3</ID>153 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>-94,-51.5</position>
<gparam>LABEL_TEXT SEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>-98,-49.5</position>
<input>
<ID>N_in2</ID>119 </input>
<input>
<ID>N_in3</ID>168 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>-95,-49.5</position>
<input>
<ID>N_in2</ID>119 </input>
<input>
<ID>N_in3</ID>167 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>-92,-49.5</position>
<input>
<ID>N_in2</ID>119 </input>
<input>
<ID>N_in3</ID>166 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>-89,-49.5</position>
<input>
<ID>N_in2</ID>119 </input>
<input>
<ID>N_in3</ID>165 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>-86,-49.5</position>
<input>
<ID>N_in2</ID>119 </input>
<input>
<ID>N_in3</ID>164 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>-83,-49.5</position>
<input>
<ID>N_in2</ID>122 </input>
<input>
<ID>N_in3</ID>163 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>GA_LED</type>
<position>-80,-49.5</position>
<input>
<ID>N_in2</ID>121 </input>
<input>
<ID>N_in3</ID>162 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>-77,-49.5</position>
<input>
<ID>N_in2</ID>120 </input>
<input>
<ID>N_in3</ID>161 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>-120,-40.5</position>
<gparam>LABEL_TEXT ADDR2MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_MUX_2x1</type>
<position>-103.5,-41</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>176 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_MUX_2x1</type>
<position>-98.5,-41</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>167 </input>
<output>
<ID>OUT</ID>175 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_MUX_2x1</type>
<position>-93.5,-41</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>174 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_MUX_2x1</type>
<position>-88.5,-41</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>165 </input>
<output>
<ID>OUT</ID>173 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_MUX_2x1</type>
<position>-83.5,-41</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>172 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_MUX_2x1</type>
<position>-78.5,-41</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>171 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_MUX_2x1</type>
<position>-73.5,-41</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>170 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_MUX_2x1</type>
<position>-68.5,-41</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>169 </output>
<input>
<ID>SEL_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-38,-173</position>
<input>
<ID>ENABLE_0</ID>57 </input>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>6 </input>
<input>
<ID>IN_4</ID>4 </input>
<input>
<ID>IN_5</ID>3 </input>
<input>
<ID>IN_6</ID>2 </input>
<input>
<ID>IN_7</ID>1 </input>
<output>
<ID>OUT_0</ID>45 </output>
<output>
<ID>OUT_1</ID>46 </output>
<output>
<ID>OUT_2</ID>47 </output>
<output>
<ID>OUT_3</ID>48 </output>
<output>
<ID>OUT_4</ID>49 </output>
<output>
<ID>OUT_5</ID>50 </output>
<output>
<ID>OUT_6</ID>51 </output>
<output>
<ID>OUT_7</ID>52 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>174</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-94.5,-31.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>19 </input>
<input>
<ID>IN_B_0</ID>169 </input>
<input>
<ID>IN_B_1</ID>170 </input>
<input>
<ID>IN_B_2</ID>171 </input>
<input>
<ID>IN_B_3</ID>172 </input>
<output>
<ID>OUT_0</ID>186 </output>
<output>
<ID>OUT_1</ID>190 </output>
<output>
<ID>OUT_2</ID>191 </output>
<output>
<ID>OUT_3</ID>189 </output>
<output>
<ID>carry_out</ID>146 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>175</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-76,-31.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>15 </input>
<input>
<ID>IN_B_0</ID>173 </input>
<input>
<ID>IN_B_1</ID>174 </input>
<input>
<ID>IN_B_2</ID>175 </input>
<input>
<ID>IN_B_3</ID>176 </input>
<output>
<ID>OUT_0</ID>192 </output>
<output>
<ID>OUT_1</ID>193 </output>
<output>
<ID>OUT_2</ID>194 </output>
<output>
<ID>OUT_3</ID>195 </output>
<input>
<ID>carry_in</ID>146 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>-60,-49.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>-106,-49.5</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>-100.5,-29.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>-69,-29</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>-32.5,-21.5</position>
<gparam>LABEL_TEXT LD.PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>-33,-14.5</position>
<gparam>LABEL_TEXT GatePC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_MUX_2x1</type>
<position>-33.5,-41.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>207 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_MUX_2x1</type>
<position>-28.5,-41.5</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>208 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_MUX_2x1</type>
<position>-23.5,-41.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>191 </input>
<output>
<ID>OUT</ID>209 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_MUX_2x1</type>
<position>-18.5,-41.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>210 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_MUX_2x1</type>
<position>-13.5,-41.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>211 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_MUX_2x1</type>
<position>-8.5,-41.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>212 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_MUX_2x1</type>
<position>-3.5,-41.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>194 </input>
<output>
<ID>OUT</ID>213 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_MUX_2x1</type>
<position>1.5,-41.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>214 </output>
<input>
<ID>SEL_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>-38.5,-45.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>4.5,-46.5</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>AE_FULLADDER_4BIT</type>
<position>8,-22</position>
<input>
<ID>IN_B_0</ID>20 </input>
<input>
<ID>IN_B_1</ID>13 </input>
<input>
<ID>IN_B_2</ID>14 </input>
<input>
<ID>IN_B_3</ID>15 </input>
<output>
<ID>OUT_0</ID>203 </output>
<output>
<ID>OUT_1</ID>204 </output>
<output>
<ID>OUT_2</ID>205 </output>
<output>
<ID>OUT_3</ID>206 </output>
<input>
<ID>carry_in</ID>197 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_FULLADDER_4BIT</type>
<position>26.5,-22</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_B_0</ID>16 </input>
<input>
<ID>IN_B_1</ID>17 </input>
<input>
<ID>IN_B_2</ID>18 </input>
<input>
<ID>IN_B_3</ID>19 </input>
<output>
<ID>OUT_0</ID>199 </output>
<output>
<ID>OUT_1</ID>200 </output>
<output>
<ID>OUT_2</ID>201 </output>
<output>
<ID>OUT_3</ID>202 </output>
<output>
<ID>carry_out</ID>197 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>5.5,-21</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>30.5,-21</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-91,-15</position>
<input>
<ID>ENABLE_0</ID>217 </input>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>194 </input>
<input>
<ID>IN_2</ID>193 </input>
<input>
<ID>IN_3</ID>192 </input>
<input>
<ID>IN_4</ID>189 </input>
<input>
<ID>IN_5</ID>191 </input>
<input>
<ID>IN_6</ID>190 </input>
<input>
<ID>IN_7</ID>186 </input>
<output>
<ID>OUT_0</ID>84 </output>
<output>
<ID>OUT_1</ID>93 </output>
<output>
<ID>OUT_2</ID>94 </output>
<output>
<ID>OUT_3</ID>95 </output>
<output>
<ID>OUT_4</ID>96 </output>
<output>
<ID>OUT_5</ID>97 </output>
<output>
<ID>OUT_6</ID>98 </output>
<output>
<ID>OUT_7</ID>99 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>-106,-14.5</position>
<gparam>LABEL_TEXT GateMAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>EE_VDD</type>
<position>117.5,8</position>
<output>
<ID>OUT_0</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>222</ID>
<type>EE_VDD</type>
<position>117.5,-7</position>
<output>
<ID>OUT_0</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>225</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>167.5,1.5</position>
<input>
<ID>ENABLE_0</ID>419 </input>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>306 </input>
<input>
<ID>IN_2</ID>301 </input>
<input>
<ID>IN_3</ID>296 </input>
<input>
<ID>IN_4</ID>291 </input>
<input>
<ID>IN_5</ID>286 </input>
<input>
<ID>IN_6</ID>279 </input>
<input>
<ID>IN_7</ID>278 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>98 </output>
<output>
<ID>OUT_2</ID>97 </output>
<output>
<ID>OUT_3</ID>96 </output>
<output>
<ID>OUT_4</ID>95 </output>
<output>
<ID>OUT_5</ID>94 </output>
<output>
<ID>OUT_6</ID>93 </output>
<output>
<ID>OUT_7</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>226</ID>
<type>GA_LED</type>
<position>81,31.5</position>
<input>
<ID>N_in0</ID>117 </input>
<input>
<ID>N_in1</ID>404 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>GA_LED</type>
<position>81,27.5</position>
<input>
<ID>N_in0</ID>118 </input>
<input>
<ID>N_in1</ID>405 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>229</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>93.5,1</position>
<input>
<ID>ENABLE_0</ID>228 </input>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>84 </input>
<output>
<ID>OUT_0</ID>236 </output>
<output>
<ID>OUT_1</ID>233 </output>
<output>
<ID>OUT_2</ID>235 </output>
<output>
<ID>OUT_3</ID>234 </output>
<output>
<ID>OUT_4</ID>238 </output>
<output>
<ID>OUT_5</ID>239 </output>
<output>
<ID>OUT_6</ID>237 </output>
<output>
<ID>OUT_7</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>230</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>93.5,-14</position>
<input>
<ID>ENABLE_0</ID>227 </input>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>84 </input>
<output>
<ID>OUT_0</ID>240 </output>
<output>
<ID>OUT_1</ID>242 </output>
<output>
<ID>OUT_2</ID>241 </output>
<output>
<ID>OUT_3</ID>243 </output>
<output>
<ID>OUT_4</ID>244 </output>
<output>
<ID>OUT_5</ID>245 </output>
<output>
<ID>OUT_6</ID>247 </output>
<output>
<ID>OUT_7</ID>246 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>231</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>93.5,-29</position>
<input>
<ID>ENABLE_0</ID>226 </input>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>84 </input>
<output>
<ID>OUT_0</ID>261 </output>
<output>
<ID>OUT_1</ID>257 </output>
<output>
<ID>OUT_2</ID>262 </output>
<output>
<ID>OUT_3</ID>260 </output>
<output>
<ID>OUT_4</ID>258 </output>
<output>
<ID>OUT_5</ID>263 </output>
<output>
<ID>OUT_6</ID>256 </output>
<output>
<ID>OUT_7</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>232</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>93.5,16</position>
<input>
<ID>ENABLE_0</ID>229 </input>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>94 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>84 </input>
<output>
<ID>OUT_0</ID>251 </output>
<output>
<ID>OUT_1</ID>248 </output>
<output>
<ID>OUT_2</ID>252 </output>
<output>
<ID>OUT_3</ID>249 </output>
<output>
<ID>OUT_4</ID>250 </output>
<output>
<ID>OUT_5</ID>253 </output>
<output>
<ID>OUT_6</ID>254 </output>
<output>
<ID>OUT_7</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>56,4.5</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>54.5,-14.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>GA_LED</type>
<position>105,31.5</position>
<input>
<ID>N_in0</ID>409 </input>
<input>
<ID>N_in1</ID>281 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>AA_LABEL</type>
<position>76,30.5</position>
<gparam>LABEL_TEXT DR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>BA_DECODER_2x4</type>
<position>87.5,31</position>
<input>
<ID>IN_0</ID>405 </input>
<input>
<ID>IN_1</ID>404 </input>
<output>
<ID>OUT_0</ID>226 </output>
<output>
<ID>OUT_1</ID>227 </output>
<output>
<ID>OUT_2</ID>228 </output>
<output>
<ID>OUT_3</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>AE_REGISTER8</type>
<position>99.5,15.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>248 </input>
<input>
<ID>IN_2</ID>252 </input>
<input>
<ID>IN_3</ID>249 </input>
<input>
<ID>IN_4</ID>250 </input>
<input>
<ID>IN_5</ID>253 </input>
<input>
<ID>IN_6</ID>254 </input>
<input>
<ID>IN_7</ID>255 </input>
<output>
<ID>OUT_0</ID>308 </output>
<output>
<ID>OUT_1</ID>302 </output>
<output>
<ID>OUT_2</ID>297 </output>
<output>
<ID>OUT_3</ID>292 </output>
<output>
<ID>OUT_4</ID>287 </output>
<output>
<ID>OUT_5</ID>282 </output>
<output>
<ID>OUT_6</ID>274 </output>
<output>
<ID>OUT_7</ID>270 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>268 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_REGISTER8</type>
<position>99.5,0.5</position>
<input>
<ID>IN_0</ID>236 </input>
<input>
<ID>IN_1</ID>233 </input>
<input>
<ID>IN_2</ID>235 </input>
<input>
<ID>IN_3</ID>234 </input>
<input>
<ID>IN_4</ID>238 </input>
<input>
<ID>IN_5</ID>239 </input>
<input>
<ID>IN_6</ID>237 </input>
<input>
<ID>IN_7</ID>232 </input>
<output>
<ID>OUT_0</ID>309 </output>
<output>
<ID>OUT_1</ID>303 </output>
<output>
<ID>OUT_2</ID>298 </output>
<output>
<ID>OUT_3</ID>293 </output>
<output>
<ID>OUT_4</ID>288 </output>
<output>
<ID>OUT_5</ID>283 </output>
<output>
<ID>OUT_6</ID>275 </output>
<output>
<ID>OUT_7</ID>271 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>267 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_REGISTER8</type>
<position>99.5,-14.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>242 </input>
<input>
<ID>IN_2</ID>241 </input>
<input>
<ID>IN_3</ID>243 </input>
<input>
<ID>IN_4</ID>244 </input>
<input>
<ID>IN_5</ID>245 </input>
<input>
<ID>IN_6</ID>247 </input>
<input>
<ID>IN_7</ID>246 </input>
<output>
<ID>OUT_0</ID>310 </output>
<output>
<ID>OUT_1</ID>304 </output>
<output>
<ID>OUT_2</ID>299 </output>
<output>
<ID>OUT_3</ID>294 </output>
<output>
<ID>OUT_4</ID>289 </output>
<output>
<ID>OUT_5</ID>284 </output>
<output>
<ID>OUT_6</ID>276 </output>
<output>
<ID>OUT_7</ID>272 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>266 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_REGISTER8</type>
<position>99.5,-29.5</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>257 </input>
<input>
<ID>IN_2</ID>262 </input>
<input>
<ID>IN_3</ID>260 </input>
<input>
<ID>IN_4</ID>258 </input>
<input>
<ID>IN_5</ID>263 </input>
<input>
<ID>IN_6</ID>256 </input>
<input>
<ID>IN_7</ID>259 </input>
<output>
<ID>OUT_0</ID>311 </output>
<output>
<ID>OUT_1</ID>305 </output>
<output>
<ID>OUT_2</ID>300 </output>
<output>
<ID>OUT_3</ID>295 </output>
<output>
<ID>OUT_4</ID>290 </output>
<output>
<ID>OUT_5</ID>285 </output>
<output>
<ID>OUT_6</ID>277 </output>
<output>
<ID>OUT_7</ID>273 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>265 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>243</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>93.5,31</position>
<input>
<ID>ENABLE_0</ID>264 </input>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>227 </input>
<input>
<ID>IN_2</ID>228 </input>
<input>
<ID>IN_3</ID>229 </input>
<output>
<ID>OUT_0</ID>265 </output>
<output>
<ID>OUT_1</ID>266 </output>
<output>
<ID>OUT_2</ID>267 </output>
<output>
<ID>OUT_3</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>244</ID>
<type>GA_LED</type>
<position>105,28.5</position>
<input>
<ID>N_in0</ID>414 </input>
<input>
<ID>N_in1</ID>280 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AE_REGISTER8</type>
<position>118.5,1</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>306 </input>
<input>
<ID>IN_2</ID>301 </input>
<input>
<ID>IN_3</ID>296 </input>
<input>
<ID>IN_4</ID>291 </input>
<input>
<ID>IN_5</ID>286 </input>
<input>
<ID>IN_6</ID>279 </input>
<input>
<ID>IN_7</ID>278 </input>
<output>
<ID>OUT_0</ID>328 </output>
<output>
<ID>OUT_1</ID>329 </output>
<output>
<ID>OUT_2</ID>330 </output>
<output>
<ID>OUT_3</ID>331 </output>
<output>
<ID>OUT_4</ID>332 </output>
<output>
<ID>OUT_5</ID>333 </output>
<output>
<ID>OUT_6</ID>334 </output>
<output>
<ID>OUT_7</ID>335 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>230 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>247</ID>
<type>AE_REGISTER8</type>
<position>118.5,-14</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>320 </input>
<input>
<ID>IN_2</ID>319 </input>
<input>
<ID>IN_3</ID>318 </input>
<input>
<ID>IN_4</ID>317 </input>
<input>
<ID>IN_5</ID>316 </input>
<input>
<ID>IN_6</ID>315 </input>
<input>
<ID>IN_7</ID>314 </input>
<output>
<ID>OUT_0</ID>324 </output>
<output>
<ID>OUT_1</ID>325 </output>
<output>
<ID>OUT_2</ID>326 </output>
<output>
<ID>OUT_3</ID>327 </output>
<output>
<ID>OUT_4</ID>339 </output>
<output>
<ID>OUT_5</ID>338 </output>
<output>
<ID>OUT_6</ID>337 </output>
<output>
<ID>OUT_7</ID>336 </output>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>load</ID>231 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>248</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>272 </input>
<input>
<ID>IN_2</ID>271 </input>
<input>
<ID>IN_3</ID>270 </input>
<output>
<ID>OUT</ID>278 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>249</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_2</ID>275 </input>
<input>
<ID>IN_3</ID>274 </input>
<output>
<ID>OUT</ID>279 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>106.5,26.5</position>
<gparam>LABEL_TEXT SR1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>285 </input>
<input>
<ID>IN_1</ID>284 </input>
<input>
<ID>IN_2</ID>283 </input>
<input>
<ID>IN_3</ID>282 </input>
<output>
<ID>OUT</ID>286 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>290 </input>
<input>
<ID>IN_1</ID>289 </input>
<input>
<ID>IN_2</ID>288 </input>
<input>
<ID>IN_3</ID>287 </input>
<output>
<ID>OUT</ID>291 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>255</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>295 </input>
<input>
<ID>IN_1</ID>294 </input>
<input>
<ID>IN_2</ID>293 </input>
<input>
<ID>IN_3</ID>292 </input>
<output>
<ID>OUT</ID>296 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>256</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>299 </input>
<input>
<ID>IN_2</ID>298 </input>
<input>
<ID>IN_3</ID>297 </input>
<output>
<ID>OUT</ID>301 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>257</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>304 </input>
<input>
<ID>IN_2</ID>303 </input>
<input>
<ID>IN_3</ID>302 </input>
<output>
<ID>OUT</ID>306 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>258</ID>
<type>AE_MUX_4x1</type>
<position>108.5,1</position>
<input>
<ID>IN_0</ID>311 </input>
<input>
<ID>IN_1</ID>310 </input>
<input>
<ID>IN_2</ID>309 </input>
<input>
<ID>IN_3</ID>308 </input>
<output>
<ID>OUT</ID>307 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>259</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>272 </input>
<input>
<ID>IN_2</ID>271 </input>
<input>
<ID>IN_3</ID>270 </input>
<output>
<ID>OUT</ID>314 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>113,26.5</position>
<gparam>LABEL_TEXT SR2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>276 </input>
<input>
<ID>IN_2</ID>275 </input>
<input>
<ID>IN_3</ID>274 </input>
<output>
<ID>OUT</ID>315 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>264</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>285 </input>
<input>
<ID>IN_1</ID>284 </input>
<input>
<ID>IN_2</ID>283 </input>
<input>
<ID>IN_3</ID>282 </input>
<output>
<ID>OUT</ID>316 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>265</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>290 </input>
<input>
<ID>IN_1</ID>289 </input>
<input>
<ID>IN_2</ID>288 </input>
<input>
<ID>IN_3</ID>287 </input>
<output>
<ID>OUT</ID>317 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>266</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>295 </input>
<input>
<ID>IN_1</ID>294 </input>
<input>
<ID>IN_2</ID>293 </input>
<input>
<ID>IN_3</ID>292 </input>
<output>
<ID>OUT</ID>318 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>267</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>299 </input>
<input>
<ID>IN_2</ID>298 </input>
<input>
<ID>IN_3</ID>297 </input>
<output>
<ID>OUT</ID>319 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>268</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>304 </input>
<input>
<ID>IN_2</ID>303 </input>
<input>
<ID>IN_3</ID>302 </input>
<output>
<ID>OUT</ID>320 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_MUX_4x1</type>
<position>108.5,-14</position>
<input>
<ID>IN_0</ID>311 </input>
<input>
<ID>IN_1</ID>310 </input>
<input>
<ID>IN_2</ID>309 </input>
<input>
<ID>IN_3</ID>308 </input>
<output>
<ID>OUT</ID>321 </output>
<input>
<ID>SEL_0</ID>313 </input>
<input>
<ID>SEL_1</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>180.5,-161</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>168.5,-160.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>AA_LABEL</type>
<position>-45,-41</position>
<gparam>LABEL_TEXT PCMUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>EE_VDD</type>
<position>36.5,-69.5</position>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>274</ID>
<type>EE_VDD</type>
<position>36.5,-89</position>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>275</ID>
<type>EE_VDD</type>
<position>36,-109</position>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>276</ID>
<type>EE_VDD</type>
<position>36.5,-128.5</position>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>277</ID>
<type>EE_VDD</type>
<position>60.5,-88.5</position>
<output>
<ID>OUT_0</ID>152 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>278</ID>
<type>EE_VDD</type>
<position>60.5,-109</position>
<output>
<ID>OUT_0</ID>177 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>279</ID>
<type>GA_LED</type>
<position>112,31.5</position>
<input>
<ID>N_in0</ID>312 </input>
<input>
<ID>N_in1</ID>121 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>GA_LED</type>
<position>112,28.5</position>
<input>
<ID>N_in0</ID>313 </input>
<input>
<ID>N_in1</ID>120 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>AA_LABEL</type>
<position>93.5,39</position>
<gparam>LABEL_TEXT LD.REG</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>287</ID>
<type>AA_LABEL</type>
<position>120,28.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>AA_LABEL</type>
<position>119.5,31.5</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>119,-23</position>
<gparam>LABEL_TEXT SR2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>AA_LABEL</type>
<position>119,11.5</position>
<gparam>LABEL_TEXT SR1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>87.5,-28</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>88,16.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>88,-1.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>88,-13</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>BA_ROM_4x4</type>
<position>54.5,-88</position>
<input>
<ID>ADDRESS_0</ID>66 </input>
<input>
<ID>ADDRESS_1</ID>61 </input>
<input>
<ID>ADDRESS_2</ID>60 </input>
<input>
<ID>ADDRESS_3</ID>59 </input>
<output>
<ID>DATA_OUT_0</ID>216 </output>
<output>
<ID>DATA_OUT_1</ID>219 </output>
<output>
<ID>DATA_OUT_2</ID>221 </output>
<output>
<ID>DATA_OUT_3</ID>218 </output>
<input>
<ID>ENABLE_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 8</lparam>
<lparam>Address:1 8</lparam>
<lparam>Address:5 6</lparam>
<lparam>Address:9 8</lparam>
<lparam>Address:10 6</lparam>
<lparam>Address:14 5</lparam></gate>
<gate>
<ID>296</ID>
<type>BA_ROM_4x4</type>
<position>54.5,-108.5</position>
<input>
<ID>ADDRESS_0</ID>66 </input>
<input>
<ID>ADDRESS_1</ID>61 </input>
<input>
<ID>ADDRESS_2</ID>60 </input>
<input>
<ID>ADDRESS_3</ID>59 </input>
<output>
<ID>DATA_OUT_0</ID>223 </output>
<output>
<ID>DATA_OUT_1</ID>322 </output>
<output>
<ID>DATA_OUT_2</ID>383 </output>
<output>
<ID>DATA_OUT_3</ID>269 </output>
<input>
<ID>ENABLE_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:1 8</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:9 8</lparam>
<lparam>Address:11 4</lparam>
<lparam>Address:14 1</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_LABEL</type>
<position>121,-119</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>305</ID>
<type>AA_LABEL</type>
<position>102,35</position>
<gparam>LABEL_TEXT ST BIT</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>AA_MUX_2x1</type>
<position>102,31.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>413 </input>
<output>
<ID>OUT</ID>409 </output>
<input>
<ID>SEL_0</ID>411 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>FF_GND</type>
<position>99,32.5</position>
<output>
<ID>OUT_0</ID>413 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_MUX_2x1</type>
<position>102,27</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>414 </output>
<input>
<ID>SEL_0</ID>411 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_LABEL</type>
<position>147,-119</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>319</ID>
<type>AE_FULLADDER_4BIT</type>
<position>151,-98</position>
<input>
<ID>IN_0</ID>328 </input>
<input>
<ID>IN_1</ID>329 </input>
<input>
<ID>IN_2</ID>330 </input>
<input>
<ID>IN_3</ID>331 </input>
<input>
<ID>IN_B_0</ID>324 </input>
<input>
<ID>IN_B_1</ID>325 </input>
<input>
<ID>IN_B_2</ID>326 </input>
<input>
<ID>IN_B_3</ID>327 </input>
<output>
<ID>OUT_0</ID>340 </output>
<output>
<ID>OUT_1</ID>341 </output>
<output>
<ID>OUT_2</ID>342 </output>
<output>
<ID>OUT_3</ID>343 </output>
<output>
<ID>carry_out</ID>323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>320</ID>
<type>AE_FULLADDER_4BIT</type>
<position>135,-98</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>333 </input>
<input>
<ID>IN_2</ID>334 </input>
<input>
<ID>IN_3</ID>335 </input>
<input>
<ID>IN_B_0</ID>339 </input>
<input>
<ID>IN_B_1</ID>338 </input>
<input>
<ID>IN_B_2</ID>337 </input>
<input>
<ID>IN_B_3</ID>336 </input>
<output>
<ID>OUT_0</ID>344 </output>
<output>
<ID>OUT_1</ID>345 </output>
<output>
<ID>OUT_2</ID>346 </output>
<output>
<ID>OUT_3</ID>347 </output>
<input>
<ID>carry_in</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>321</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>143,-106</position>
<input>
<ID>ENABLE_0</ID>372 </input>
<input>
<ID>IN_0</ID>347 </input>
<input>
<ID>IN_1</ID>346 </input>
<input>
<ID>IN_2</ID>345 </input>
<input>
<ID>IN_3</ID>344 </input>
<input>
<ID>IN_4</ID>343 </input>
<input>
<ID>IN_5</ID>342 </input>
<input>
<ID>IN_6</ID>341 </input>
<input>
<ID>IN_7</ID>340 </input>
<output>
<ID>OUT_0</ID>356 </output>
<output>
<ID>OUT_1</ID>357 </output>
<output>
<ID>OUT_2</ID>358 </output>
<output>
<ID>OUT_3</ID>359 </output>
<output>
<ID>OUT_4</ID>360 </output>
<output>
<ID>OUT_5</ID>361 </output>
<output>
<ID>OUT_6</ID>362 </output>
<output>
<ID>OUT_7</ID>363 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>322</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>337 </input>
<input>
<ID>IN_1</ID>334 </input>
<output>
<ID>OUT</ID>349 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>336 </input>
<input>
<ID>IN_1</ID>335 </input>
<output>
<ID>OUT</ID>348 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>116,-106</position>
<input>
<ID>ENABLE_0</ID>374 </input>
<input>
<ID>IN_0</ID>348 </input>
<input>
<ID>IN_1</ID>349 </input>
<input>
<ID>IN_2</ID>350 </input>
<input>
<ID>IN_3</ID>351 </input>
<input>
<ID>IN_4</ID>352 </input>
<input>
<ID>IN_5</ID>353 </input>
<input>
<ID>IN_6</ID>354 </input>
<input>
<ID>IN_7</ID>355 </input>
<output>
<ID>OUT_0</ID>356 </output>
<output>
<ID>OUT_1</ID>357 </output>
<output>
<ID>OUT_2</ID>358 </output>
<output>
<ID>OUT_3</ID>359 </output>
<output>
<ID>OUT_4</ID>360 </output>
<output>
<ID>OUT_5</ID>361 </output>
<output>
<ID>OUT_6</ID>362 </output>
<output>
<ID>OUT_7</ID>363 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>338 </input>
<input>
<ID>IN_1</ID>333 </input>
<output>
<ID>OUT</ID>350 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>326</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>339 </input>
<input>
<ID>IN_1</ID>332 </input>
<output>
<ID>OUT</ID>351 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>327 </input>
<input>
<ID>IN_1</ID>331 </input>
<output>
<ID>OUT</ID>352 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>353 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>325 </input>
<input>
<ID>IN_1</ID>329 </input>
<output>
<ID>OUT</ID>354 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AA_AND2</type>
<position>116,-98</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>355 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>134,-110</position>
<input>
<ID>ENABLE_0</ID>373 </input>
<input>
<ID>IN_0</ID>356 </input>
<input>
<ID>IN_1</ID>357 </input>
<input>
<ID>IN_2</ID>358 </input>
<input>
<ID>IN_3</ID>359 </input>
<input>
<ID>IN_4</ID>360 </input>
<input>
<ID>IN_5</ID>361 </input>
<input>
<ID>IN_6</ID>362 </input>
<input>
<ID>IN_7</ID>363 </input>
<output>
<ID>OUT_0</ID>364 </output>
<output>
<ID>OUT_1</ID>365 </output>
<output>
<ID>OUT_2</ID>366 </output>
<output>
<ID>OUT_3</ID>367 </output>
<output>
<ID>OUT_4</ID>368 </output>
<output>
<ID>OUT_5</ID>369 </output>
<output>
<ID>OUT_6</ID>370 </output>
<output>
<ID>OUT_7</ID>371 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>333</ID>
<type>GA_LED</type>
<position>123.5,-114</position>
<input>
<ID>N_in2</ID>84 </input>
<input>
<ID>N_in3</ID>364 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>334</ID>
<type>GA_LED</type>
<position>126.5,-114</position>
<input>
<ID>N_in2</ID>93 </input>
<input>
<ID>N_in3</ID>365 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>335</ID>
<type>GA_LED</type>
<position>129.5,-114</position>
<input>
<ID>N_in2</ID>94 </input>
<input>
<ID>N_in3</ID>366 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>336</ID>
<type>GA_LED</type>
<position>132.5,-114</position>
<input>
<ID>N_in2</ID>95 </input>
<input>
<ID>N_in3</ID>367 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>337</ID>
<type>GA_LED</type>
<position>135.5,-114</position>
<input>
<ID>N_in2</ID>96 </input>
<input>
<ID>N_in3</ID>368 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>GA_LED</type>
<position>138.5,-114</position>
<input>
<ID>N_in2</ID>97 </input>
<input>
<ID>N_in3</ID>369 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>339</ID>
<type>GA_LED</type>
<position>141.5,-114</position>
<input>
<ID>N_in2</ID>98 </input>
<input>
<ID>N_in3</ID>370 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>340</ID>
<type>GA_LED</type>
<position>144.5,-114</position>
<input>
<ID>N_in2</ID>99 </input>
<input>
<ID>N_in3</ID>371 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>AE_SMALL_INVERTER</type>
<position>123,-106</position>
<input>
<ID>IN_0</ID>372 </input>
<output>
<ID>OUT_0</ID>374 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_AND2</type>
<position>-13.5,-99</position>
<input>
<ID>IN_0</ID>377 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>375 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_LABEL</type>
<position>-49.5,-43.5</position>
<gparam>LABEL_TEXT OFF = +1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>EE_VDD</type>
<position>24.5,-13</position>
<output>
<ID>OUT_0</ID>378 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>348</ID>
<type>AA_LABEL</type>
<position>-118,-44</position>
<gparam>LABEL_TEXT OFF = SEXT3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>AA_LABEL</type>
<position>167.5,-86</position>
<gparam>LABEL_TEXT On =ADD</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>350</ID>
<type>AA_LABEL</type>
<position>151,-109.5</position>
<gparam>LABEL_TEXT GateALU</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>355</ID>
<type>AA_LABEL</type>
<position>137.5,12</position>
<gparam>LABEL_TEXT SRC-Mem Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AA_LABEL</type>
<position>30.5,-125</position>
<gparam>LABEL_TEXT ROM4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>357</ID>
<type>AA_LABEL</type>
<position>30.5,-106</position>
<gparam>LABEL_TEXT ROM3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>358</ID>
<type>AA_LABEL</type>
<position>55.5,-85</position>
<gparam>LABEL_TEXT ROM5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>359</ID>
<type>AA_LABEL</type>
<position>55,-105.5</position>
<gparam>LABEL_TEXT ROM6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>362</ID>
<type>AA_AND2</type>
<position>-104.5,-143</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>BB_CLOCK</type>
<position>-111.5,-142</position>
<output>
<ID>CLK</ID>380 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>366</ID>
<type>AA_TOGGLE</type>
<position>-111,-148.5</position>
<output>
<ID>OUT_0</ID>381 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,-181.5,-6.5,-181.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_7</name></connection>
<intersection>-41.5 6</intersection>
<intersection>-14 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-41.5,-181.5,-41.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_7</name></connection>
<intersection>-181.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-14,-182,-14,-181.5</points>
<connection>
<GID>73</GID>
<name>OUT_7</name></connection>
<intersection>-181.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40.5,-182.5,-6.5,-182.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_6</name></connection>
<intersection>-40.5 4</intersection>
<intersection>-14 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-40.5,-182.5,-40.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_6</name></connection>
<intersection>-182.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-14,-183,-14,-182.5</points>
<connection>
<GID>73</GID>
<name>OUT_6</name></connection>
<intersection>-182.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39.5,-183.5,-6.5,-183.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_5</name></connection>
<intersection>-39.5 2</intersection>
<intersection>-14 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-39.5,-183.5,-39.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_5</name></connection>
<intersection>-183.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-14,-184,-14,-183.5</points>
<connection>
<GID>73</GID>
<name>OUT_5</name></connection>
<intersection>-183.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38.5,-184.5,-6.5,-184.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_4</name></connection>
<intersection>-38.5 4</intersection>
<intersection>-14 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-38.5,-184.5,-38.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_4</name></connection>
<intersection>-184.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-14,-185,-14,-184.5</points>
<connection>
<GID>73</GID>
<name>OUT_4</name></connection>
<intersection>-184.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.38498e-008,-118.5,-2.38498e-008,-116.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-116.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>2,-116.5,2,-114.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>-116.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2.38498e-008,-116.5,2,-116.5</points>
<intersection>-2.38498e-008 0</intersection>
<intersection>2 1</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-166,-44.5,-104</points>
<intersection>-166 5</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,-104,53.5,-104</points>
<intersection>-44.5 0</intersection>
<intersection>53.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>53.5,-104,53.5,-103</points>
<intersection>-104 1</intersection>
<intersection>-103 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>53.5,-103,55,-103</points>
<intersection>53.5 2</intersection>
<intersection>55 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>55,-103,55,-102</points>
<connection>
<GID>138</GID>
<name>OUT_2</name></connection>
<intersection>-103 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-44.5,-166,-43.5,-166</points>
<connection>
<GID>11</GID>
<name>load</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-118.5,2,-118.5</points>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37.5,-185.5,-6.5,-185.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_3</name></connection>
<intersection>-37.5 4</intersection>
<intersection>-14 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-37.5,-185.5,-37.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_3</name></connection>
<intersection>-185.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-14,-186,-14,-185.5</points>
<connection>
<GID>73</GID>
<name>OUT_3</name></connection>
<intersection>-185.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-118.5,9.5,-118.5</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-186.5,-6.5,-186.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_2</name></connection>
<intersection>-36.5 4</intersection>
<intersection>-14 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-36.5,-186.5,-36.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_2</name></connection>
<intersection>-186.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-14,-187,-14,-186.5</points>
<connection>
<GID>73</GID>
<name>OUT_2</name></connection>
<intersection>-186.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35.5,-187.5,-6.5,-187.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_1</name></connection>
<intersection>-35.5 4</intersection>
<intersection>-14 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-35.5,-187.5,-35.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>-187.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-14,-188,-14,-187.5</points>
<connection>
<GID>73</GID>
<name>OUT_1</name></connection>
<intersection>-187.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-34.5,-188.5,-6.5,-188.5</points>
<connection>
<GID>52</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>DATA_IN_0</name></connection>
<intersection>-34.5 4</intersection>
<intersection>-14 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-34.5,-188.5,-34.5,-175</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-14,-189,-14,-188.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-188.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-180,-3,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_0</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-169,-2.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-3 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80.5,-194.5,-80.5,-167</points>
<intersection>-194.5 19</intersection>
<intersection>-179.5 1</intersection>
<intersection>-167 26</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-89.5,-179.5,-30,-179.5</points>
<intersection>-89.5 5</intersection>
<intersection>-80.5 0</intersection>
<intersection>-30 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-30,-179.5,-30,-145</points>
<intersection>-179.5 1</intersection>
<intersection>-164 77</intersection>
<intersection>-145 12</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-89.5,-179.5,-89.5,-143</points>
<intersection>-179.5 1</intersection>
<intersection>-167 26</intersection>
<intersection>-143 25</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-30,-145,-25,-145</points>
<connection>
<GID>56</GID>
<name>clock</name></connection>
<intersection>-30 4</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-80.5,-194.5,101,-194.5</points>
<intersection>-80.5 0</intersection>
<intersection>2 20</intersection>
<intersection>101 40</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>2,-194.5,2,-190</points>
<connection>
<GID>52</GID>
<name>write_clock</name></connection>
<intersection>-194.5 19</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>-101.5,-143,-89.5,-143</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<intersection>-89.5 5</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-89.5,-167,-32.5,-167</points>
<intersection>-89.5 5</intersection>
<intersection>-80.5 0</intersection>
<intersection>-57 34</intersection>
<intersection>-32.5 78</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-57.5,-88,-29,-88</points>
<intersection>-57.5 62</intersection>
<intersection>-57 34</intersection>
<intersection>-42.5 63</intersection>
<intersection>-29 64</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>-57,-167,-57,-88</points>
<intersection>-167 26</intersection>
<intersection>-88 28</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>101,-194.5,101,-38.5</points>
<intersection>-194.5 19</intersection>
<intersection>-38.5 45</intersection></vsegment>
<vsegment>
<ID>41</ID>
<points>95.5,-38.5,95.5,10.5</points>
<intersection>-38.5 45</intersection>
<intersection>-34.5 42</intersection>
<intersection>-19.5 55</intersection>
<intersection>-4.5 47</intersection>
<intersection>10.5 49</intersection></vsegment>
<hsegment>
<ID>42</ID>
<points>95.5,-34.5,98.5,-34.5</points>
<connection>
<GID>242</GID>
<name>clock</name></connection>
<intersection>95.5 41</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>95.5,-38.5,112.5,-38.5</points>
<intersection>95.5 41</intersection>
<intersection>101 40</intersection>
<intersection>112.5 53</intersection></hsegment>
<hsegment>
<ID>47</ID>
<points>95.5,-4.5,98.5,-4.5</points>
<connection>
<GID>240</GID>
<name>clock</name></connection>
<intersection>95.5 41</intersection></hsegment>
<hsegment>
<ID>49</ID>
<points>95.5,10.5,98.5,10.5</points>
<connection>
<GID>239</GID>
<name>clock</name></connection>
<intersection>95.5 41</intersection></hsegment>
<vsegment>
<ID>53</ID>
<points>112.5,-38.5,112.5,-19</points>
<intersection>-38.5 45</intersection>
<intersection>-19 58</intersection></vsegment>
<hsegment>
<ID>55</ID>
<points>95.5,-19.5,98.5,-19.5</points>
<connection>
<GID>241</GID>
<name>clock</name></connection>
<intersection>95.5 41</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>112.5,-19,117.5,-19</points>
<connection>
<GID>247</GID>
<name>clock</name></connection>
<intersection>112.5 53</intersection>
<intersection>117.5 81</intersection></hsegment>
<vsegment>
<ID>62</ID>
<points>-57.5,-88,-57.5,-81</points>
<connection>
<GID>102</GID>
<name>clock</name></connection>
<intersection>-88 28</intersection></vsegment>
<vsegment>
<ID>63</ID>
<points>-42.5,-88,-42.5,-81</points>
<connection>
<GID>112</GID>
<name>clock</name></connection>
<intersection>-88 28</intersection></vsegment>
<vsegment>
<ID>64</ID>
<points>-29,-88,-29,-78.5</points>
<connection>
<GID>114</GID>
<name>clock</name></connection>
<intersection>-88 28</intersection>
<intersection>-78.5 70</intersection></vsegment>
<hsegment>
<ID>70</ID>
<points>-29,-78.5,26,-78.5</points>
<connection>
<GID>121</GID>
<name>clock</name></connection>
<intersection>-29 64</intersection>
<intersection>-16 82</intersection>
<intersection>26 71</intersection></hsegment>
<vsegment>
<ID>71</ID>
<points>26,-137,26,-78.5</points>
<connection>
<GID>124</GID>
<name>clock</name></connection>
<connection>
<GID>135</GID>
<name>clock</name></connection>
<intersection>-117 72</intersection>
<intersection>-97 74</intersection>
<intersection>-78.5 70</intersection></vsegment>
<hsegment>
<ID>72</ID>
<points>25.5,-117,26,-117</points>
<connection>
<GID>132</GID>
<name>clock</name></connection>
<intersection>26 71</intersection></hsegment>
<hsegment>
<ID>74</ID>
<points>26,-97,50,-97</points>
<connection>
<GID>138</GID>
<name>clock</name></connection>
<intersection>26 71</intersection>
<intersection>50 75</intersection></hsegment>
<vsegment>
<ID>75</ID>
<points>50,-119,50,-97</points>
<connection>
<GID>140</GID>
<name>clock</name></connection>
<intersection>-97 74</intersection></vsegment>
<hsegment>
<ID>77</ID>
<points>-30,-164,-4.5,-164</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>-30 4</intersection></hsegment>
<vsegment>
<ID>78</ID>
<points>-32.5,-167,-32.5,-166</points>
<connection>
<GID>11</GID>
<name>clock</name></connection>
<intersection>-167 26</intersection></vsegment>
<vsegment>
<ID>81</ID>
<points>117.5,-19,117.5,-4</points>
<connection>
<GID>246</GID>
<name>clock</name></connection>
<intersection>-19 58</intersection></vsegment>
<vsegment>
<ID>82</ID>
<points>-16,-78.5,-16,-22</points>
<intersection>-78.5 70</intersection>
<intersection>-22 83</intersection></vsegment>
<hsegment>
<ID>83</ID>
<points>-16,-22,-13,-22</points>
<connection>
<GID>60</GID>
<name>clock</name></connection>
<intersection>-16 82</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-36,-22.5,-15.5</points>
<intersection>-36 3</intersection>
<intersection>-15.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-73,-36,-22.5,-36</points>
<intersection>-73 4</intersection>
<intersection>-22.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-73,-36,-73,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-22.5,-15.5,12,-15.5</points>
<intersection>-22.5 0</intersection>
<intersection>-20 8</intersection>
<intersection>12 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>12,-18,12,-15.5</points>
<connection>
<GID>198</GID>
<name>IN_B_1</name></connection>
<intersection>-15.5 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-20,-17,-20,-14</points>
<connection>
<GID>62</GID>
<name>IN_5</name></connection>
<connection>
<GID>60</GID>
<name>OUT_5</name></connection>
<intersection>-15.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-36.5,-22.5,-15.5</points>
<intersection>-36.5 3</intersection>
<intersection>-17 9</intersection>
<intersection>-15.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-72,-36.5,-22.5,-36.5</points>
<intersection>-72 4</intersection>
<intersection>-22.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-72,-36.5,-72,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_2</name></connection>
<intersection>-36.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-22.5,-15.5,11,-15.5</points>
<intersection>-22.5 0</intersection>
<intersection>-21 8</intersection>
<intersection>11 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>11,-18,11,-15.5</points>
<connection>
<GID>198</GID>
<name>IN_B_2</name></connection>
<intersection>-15.5 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-21,-15.5,-21,-14</points>
<connection>
<GID>62</GID>
<name>IN_6</name></connection>
<intersection>-15.5 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-22.5,-17,-21,-17</points>
<connection>
<GID>60</GID>
<name>OUT_6</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,30.5,83,31.5</points>
<intersection>30.5 2</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,31.5,83,31.5</points>
<connection>
<GID>226</GID>
<name>N_in1</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,30.5,84.5,30.5</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-35.5,-23,-15.5</points>
<intersection>-35.5 3</intersection>
<intersection>-17 10</intersection>
<intersection>-15.5 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-71,-35.5,-23,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_3</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-23,-15.5,10,-15.5</points>
<intersection>-23 0</intersection>
<intersection>-22 9</intersection>
<intersection>10 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>10,-18,10,-15.5</points>
<connection>
<GID>198</GID>
<name>IN_B_3</name></connection>
<intersection>-15.5 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-22,-15.5,-22,-14</points>
<connection>
<GID>62</GID>
<name>IN_7</name></connection>
<intersection>-15.5 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-23,-17,-22,-17</points>
<connection>
<GID>60</GID>
<name>OUT_7</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,27.5,83,29.5</points>
<intersection>27.5 2</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,29.5,84.5,29.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,27.5,83,27.5</points>
<connection>
<GID>227</GID>
<name>N_in1</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-36,-23,-15.5</points>
<intersection>-36 1</intersection>
<intersection>-15.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-92.5,-36,-23,-36</points>
<intersection>-92.5 2</intersection>
<intersection>-23 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-92.5,-36,-92.5,-35.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-23,-15.5,31.5,-15.5</points>
<intersection>-23 0</intersection>
<intersection>-15 6</intersection>
<intersection>31.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31.5,-18,31.5,-15.5</points>
<connection>
<GID>199</GID>
<name>IN_B_0</name></connection>
<intersection>-15.5 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-15,-17,-15,-14</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-36,-23,-15.5</points>
<intersection>-36 3</intersection>
<intersection>-15.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-91.5,-36,-23,-36</points>
<intersection>-91.5 4</intersection>
<intersection>-23 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-91.5,-36,-91.5,-35.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-23,-15.5,30.5,-15.5</points>
<intersection>-23 0</intersection>
<intersection>-16 8</intersection>
<intersection>30.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>30.5,-18,30.5,-15.5</points>
<connection>
<GID>199</GID>
<name>IN_B_1</name></connection>
<intersection>-15.5 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-16,-17,-16,-14</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<connection>
<GID>60</GID>
<name>OUT_1</name></connection>
<intersection>-15.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-36,-23,-15.5</points>
<intersection>-36 3</intersection>
<intersection>-15.5 6</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-90.5,-36,-23,-36</points>
<intersection>-90.5 4</intersection>
<intersection>-23 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-90.5,-36,-90.5,-35.5</points>
<connection>
<GID>174</GID>
<name>IN_2</name></connection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-23,-15.5,29.5,-15.5</points>
<intersection>-23 0</intersection>
<intersection>-17 8</intersection>
<intersection>29.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29.5,-18,29.5,-15.5</points>
<connection>
<GID>199</GID>
<name>IN_B_2</name></connection>
<intersection>-15.5 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-17,-17,-17,-14</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<connection>
<GID>60</GID>
<name>OUT_2</name></connection>
<intersection>-15.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-89.5,-29.5,-28,-29.5</points>
<intersection>-89.5 4</intersection>
<intersection>-28 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-89.5,-35.5,-89.5,-29.5</points>
<connection>
<GID>174</GID>
<name>IN_3</name></connection>
<intersection>-29.5 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-28,-29.5,-28,-18.5</points>
<intersection>-29.5 3</intersection>
<intersection>-18.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-28,-18.5,-18.5,-18.5</points>
<intersection>-28 8</intersection>
<intersection>-18.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-18.5,-18.5,-18.5,-17</points>
<intersection>-18.5 9</intersection>
<intersection>-17 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-18.5,-17,28.5,-17</points>
<connection>
<GID>60</GID>
<name>OUT_3</name></connection>
<intersection>-18.5 10</intersection>
<intersection>-18 13</intersection>
<intersection>28.5 14</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-18,-17,-18,-14</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>-17 11</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>28.5,-18,28.5,-17</points>
<connection>
<GID>199</GID>
<name>IN_B_3</name></connection>
<intersection>-17 11</intersection></vsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,31.5,104,31.5</points>
<connection>
<GID>235</GID>
<name>N_in0</name></connection>
<connection>
<GID>307</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-36,-22.5,-15.5</points>
<intersection>-36 1</intersection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,-36,-22.5,-36</points>
<intersection>-74 2</intersection>
<intersection>-22.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-74,-36,-74,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-22.5,-15.5,13,-15.5</points>
<intersection>-22.5 0</intersection>
<intersection>-19 6</intersection>
<intersection>13 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>13,-18,13,-15.5</points>
<connection>
<GID>198</GID>
<name>IN_B_0</name></connection>
<intersection>-15.5 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-19,-17,-19,-14</points>
<connection>
<GID>62</GID>
<name>IN_4</name></connection>
<connection>
<GID>60</GID>
<name>OUT_4</name></connection>
<intersection>-15.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36,-142.5,29,-142.5</points>
<intersection>-36 4</intersection>
<intersection>29 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-36,-145,-36,-142.5</points>
<connection>
<GID>56</GID>
<name>load</name></connection>
<intersection>-142.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>29,-142.5,29,-142</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>-142.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-102.5,97,34</points>
<intersection>-102.5 2</intersection>
<intersection>34 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31,-102.5,97,-102.5</points>
<connection>
<GID>124</GID>
<name>OUT_2</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>97,34,102,34</points>
<connection>
<GID>307</GID>
<name>SEL_0</name></connection>
<intersection>97 0</intersection>
<intersection>102 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,29.5,102,34</points>
<connection>
<GID>316</GID>
<name>SEL_0</name></connection>
<intersection>34 3</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-142,32,-24.5</points>
<connection>
<GID>135</GID>
<name>OUT_3</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-24.5,32,-24.5</points>
<intersection>-24 4</intersection>
<intersection>32 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-24,-24.5,-24,-22</points>
<connection>
<GID>60</GID>
<name>load</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-123,40.5,-8</points>
<intersection>-123 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-123,40.5,-123</points>
<intersection>30.5 11</intersection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-8,40.5,-8</points>
<intersection>-23.5 4</intersection>
<intersection>40.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-23.5,-12,-23.5,-8</points>
<connection>
<GID>62</GID>
<name>ENABLE_0</name></connection>
<intersection>-8 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>30.5,-123,30.5,-122</points>
<connection>
<GID>132</GID>
<name>OUT_2</name></connection>
<intersection>-123 1</intersection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,32.5,100,32.5</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,27,104,28.5</points>
<connection>
<GID>244</GID>
<name>N_in0</name></connection>
<connection>
<GID>316</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-180,4,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_7</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-169,4.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_7</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-180,3,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_6</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-169,3.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_6</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-180,2,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_5</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-169,2.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_5</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-180,1,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_4</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-169,1.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_4</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-58,167.5,6.5</points>
<connection>
<GID>225</GID>
<name>ENABLE_0</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45.5,-122.5,45.5,-58</points>
<intersection>-122.5 3</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-58,167.5,-58</points>
<intersection>45.5 1</intersection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>45.5,-122.5,53,-122.5</points>
<intersection>45.5 1</intersection>
<intersection>53 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53,-124,53,-122.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-122.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.96046e-008,-180,-5.96046e-008,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_3</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.96046e-008,-169,0.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-5.96046e-008 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-180,-1,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_2</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-169,-0.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-180,-2,-169</points>
<connection>
<GID>52</GID>
<name>ADDRESS_1</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2,-169,-1.5,-169</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-161,-39.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_5</name></connection>
<connection>
<GID>22</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40.5,-161,-40.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_6</name></connection>
<connection>
<GID>22</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,-161,-41.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_7</name></connection>
<connection>
<GID>22</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-161,-34.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,-120.5,17,-120.5</points>
<connection>
<GID>80</GID>
<name>SEL_0</name></connection>
<connection>
<GID>77</GID>
<name>SEL_0</name></connection>
<connection>
<GID>74</GID>
<name>SEL_0</name></connection>
<connection>
<GID>78</GID>
<name>SEL_0</name></connection>
<intersection>17 29</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>17,-120.5,17,-103.5</points>
<intersection>-120.5 1</intersection>
<intersection>-103.5 30</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>17,-103.5,29,-103.5</points>
<intersection>17 29</intersection>
<intersection>29 36</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>29,-103.5,29,-102.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>-103.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-161,-35.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_1</name></connection>
<connection>
<GID>22</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-161,-36.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_2</name></connection>
<connection>
<GID>22</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37.5,-161,-37.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_3</name></connection>
<connection>
<GID>22</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38.5,-161,-38.5,-161</points>
<connection>
<GID>11</GID>
<name>OUT_4</name></connection>
<connection>
<GID>22</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-171,-34.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-171,-35.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<connection>
<GID>173</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-171,-36.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_2</name></connection>
<connection>
<GID>173</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37.5,-171,-37.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_3</name></connection>
<connection>
<GID>173</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38.5,-171,-38.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_4</name></connection>
<connection>
<GID>173</GID>
<name>OUT_4</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-171,-39.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_5</name></connection>
<connection>
<GID>173</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40.5,-171,-40.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_6</name></connection>
<connection>
<GID>173</GID>
<name>OUT_6</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,-171,-41.5,-169</points>
<connection>
<GID>11</GID>
<name>IN_7</name></connection>
<connection>
<GID>173</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-159,-43,-123</points>
<connection>
<GID>22</GID>
<name>ENABLE_0</name></connection>
<intersection>-123 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-43,-123,28.5,-123</points>
<intersection>-43 0</intersection>
<intersection>28.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>28.5,-123,28.5,-122</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>-123 3</intersection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>1,-191.5,57.5,-191.5</points>
<intersection>1 9</intersection>
<intersection>57.5 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>57.5,-191.5,57.5,-103.5</points>
<intersection>-191.5 0</intersection>
<intersection>-103.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>53,-103.5,57.5,-103.5</points>
<intersection>53 5</intersection>
<intersection>57.5 1</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53,-103.5,53,-102</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-103.5 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>1,-191.5,1,-190</points>
<connection>
<GID>52</GID>
<name>write_enable</name></connection>
<intersection>-191.5 0</intersection>
<intersection>-191 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-16,-191,1,-191</points>
<intersection>-16 13</intersection>
<intersection>1 9</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-16,-191,-16,-180.5</points>
<connection>
<GID>73</GID>
<name>ENABLE_0</name></connection>
<intersection>-191 12</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.96046e-008,-192.5,60,-192.5</points>
<intersection>5.96046e-008 4</intersection>
<intersection>60 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60,-192.5,60,-102.5</points>
<intersection>-192.5 1</intersection>
<intersection>-102.5 8</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>5.96046e-008,-192.5,5.96046e-008,-190</points>
<connection>
<GID>52</GID>
<name>ENABLE_0</name></connection>
<intersection>-192.5 1</intersection>
<intersection>-190.5 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>54,-102.5,60,-102.5</points>
<intersection>54 9</intersection>
<intersection>60 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>54,-102.5,54,-102</points>
<connection>
<GID>138</GID>
<name>OUT_1</name></connection>
<intersection>-102.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-43.5,-190.5,5.96046e-008,-190.5</points>
<intersection>-43.5 11</intersection>
<intersection>5.96046e-008 4</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-43.5,-190.5,-43.5,-173</points>
<intersection>-190.5 10</intersection>
<intersection>-173 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-43.5,-173,-43,-173</points>
<connection>
<GID>173</GID>
<name>ENABLE_0</name></connection>
<intersection>-43.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-124.5,19,-67.5</points>
<intersection>-124.5 2</intersection>
<intersection>-107 4</intersection>
<intersection>-87 11</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-67.5,25.5,-67.5</points>
<connection>
<GID>127</GID>
<name>ADDRESS_3</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-124.5,48.5,-124.5</points>
<intersection>-13.5 3</intersection>
<intersection>19 0</intersection>
<intersection>22.5 6</intersection>
<intersection>48.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-13.5,-124.5,-13.5,-122.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-107,25,-107</points>
<connection>
<GID>131</GID>
<name>ADDRESS_3</name></connection>
<intersection>19 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>22.5,-126.5,22.5,-124.5</points>
<intersection>-126.5 12</intersection>
<intersection>-124.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>48.5,-124.5,48.5,-86.5</points>
<intersection>-124.5 2</intersection>
<intersection>-107 9</intersection>
<intersection>-86.5 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>48.5,-107,49.5,-107</points>
<connection>
<GID>296</GID>
<name>ADDRESS_3</name></connection>
<intersection>48.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>48.5,-86.5,49.5,-86.5</points>
<connection>
<GID>295</GID>
<name>ADDRESS_3</name></connection>
<intersection>48.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>19,-87,25.5,-87</points>
<connection>
<GID>129</GID>
<name>ADDRESS_3</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>22.5,-126.5,25,-126.5</points>
<connection>
<GID>125</GID>
<name>ADDRESS_3</name></connection>
<intersection>22.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-127.5,20,-68.5</points>
<intersection>-127.5 5</intersection>
<intersection>-124 2</intersection>
<intersection>-108 4</intersection>
<intersection>-88 13</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-68.5,25.5,-68.5</points>
<connection>
<GID>127</GID>
<name>ADDRESS_2</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7,-124,20,-124</points>
<intersection>-7 3</intersection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-7,-124,-7,-122.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,-108,25,-108</points>
<connection>
<GID>131</GID>
<name>ADDRESS_2</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>20,-127.5,25,-127.5</points>
<connection>
<GID>125</GID>
<name>ADDRESS_2</name></connection>
<intersection>20 0</intersection>
<intersection>24.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>24.5,-132,24.5,-127.5</points>
<intersection>-132 9</intersection>
<intersection>-127.5 5</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>24.5,-132,49.5,-132</points>
<intersection>24.5 6</intersection>
<intersection>48.5 11</intersection>
<intersection>49.5 14</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>48.5,-132,48.5,-87.5</points>
<intersection>-132 9</intersection>
<intersection>-87.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>48.5,-87.5,49.5,-87.5</points>
<connection>
<GID>295</GID>
<name>ADDRESS_2</name></connection>
<intersection>48.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>20,-88,25.5,-88</points>
<connection>
<GID>129</GID>
<name>ADDRESS_2</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>49.5,-132,49.5,-108</points>
<connection>
<GID>296</GID>
<name>ADDRESS_2</name></connection>
<intersection>-132 9</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-126,20.5,-69.5</points>
<intersection>-126 5</intersection>
<intersection>-124.5 2</intersection>
<intersection>-109 4</intersection>
<intersection>-89 11</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-69.5,25.5,-69.5</points>
<connection>
<GID>127</GID>
<name>ADDRESS_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-124.5,20.5,-124.5</points>
<intersection>1 3</intersection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1,-124.5,1,-122.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20.5,-109,25,-109</points>
<connection>
<GID>131</GID>
<name>ADDRESS_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>20.5,-126,48.5,-126</points>
<intersection>20.5 0</intersection>
<intersection>23.5 10</intersection>
<intersection>48.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>48.5,-126,48.5,-88.5</points>
<intersection>-126 5</intersection>
<intersection>-109 9</intersection>
<intersection>-88.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>48.5,-88.5,49.5,-88.5</points>
<connection>
<GID>295</GID>
<name>ADDRESS_1</name></connection>
<intersection>48.5 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>48.5,-109,49.5,-109</points>
<connection>
<GID>296</GID>
<name>ADDRESS_1</name></connection>
<intersection>48.5 6</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>23.5,-128.5,23.5,-126</points>
<intersection>-128.5 12</intersection>
<intersection>-126 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>20.5,-89,25.5,-89</points>
<connection>
<GID>129</GID>
<name>ADDRESS_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>23.5,-128.5,25,-128.5</points>
<connection>
<GID>125</GID>
<name>ADDRESS_1</name></connection>
<intersection>23.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>1,-108.5,1,-84</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>1,-84,30,-84</points>
<intersection>1 1</intersection>
<intersection>30 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30,-84,30,-83.5</points>
<connection>
<GID>121</GID>
<name>OUT_1</name></connection>
<intersection>-84 2</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-129.5,21.5,-70.5</points>
<intersection>-129.5 6</intersection>
<intersection>-125 2</intersection>
<intersection>-110 4</intersection>
<intersection>-90 11</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-70.5,25.5,-70.5</points>
<connection>
<GID>127</GID>
<name>ADDRESS_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-125,21.5,-125</points>
<intersection>8.5 3</intersection>
<intersection>21.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8.5,-125,8.5,-122.5</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>-125 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-110,25,-110</points>
<connection>
<GID>131</GID>
<name>ADDRESS_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21.5,-129.5,48.5,-129.5</points>
<connection>
<GID>125</GID>
<name>ADDRESS_0</name></connection>
<intersection>21.5 0</intersection>
<intersection>48.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>48.5,-129.5,48.5,-89.5</points>
<intersection>-129.5 6</intersection>
<intersection>-110 10</intersection>
<intersection>-89.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>48.5,-89.5,49.5,-89.5</points>
<connection>
<GID>295</GID>
<name>ADDRESS_0</name></connection>
<intersection>48.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>48.5,-110,49.5,-110</points>
<connection>
<GID>296</GID>
<name>ADDRESS_0</name></connection>
<intersection>48.5 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>21.5,-90,25.5,-90</points>
<connection>
<GID>129</GID>
<name>ADDRESS_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>3,-108.5,3,-108.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-102.5,2.5,-78.5</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>-102.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>2,-102.5,2.5,-102.5</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-116.5,-12.5,-115</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-116.5,-12.5,-116.5</points>
<intersection>-14.5 7</intersection>
<intersection>-12.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-14.5,-118.5,-14.5,-116.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-116.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>7.5,-118.5,7.5,-84</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-84,29,-84</points>
<intersection>7.5 1</intersection>
<intersection>29 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>29,-84,29,-83.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>-84 2</intersection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-102.5,4,-101.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-101.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>4,-101.5,30,-101.5</points>
<intersection>4 0</intersection>
<intersection>30 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30,-102.5,30,-101.5</points>
<connection>
<GID>124</GID>
<name>OUT_1</name></connection>
<intersection>-101.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-140,-34,-118</points>
<connection>
<GID>56</GID>
<name>OUT_7</name></connection>
<intersection>-118 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-34,-118,-12.5,-118</points>
<intersection>-34 0</intersection>
<intersection>-12.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-12.5,-118.5,-12.5,-118</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>-118 3</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-140,-33,-117</points>
<connection>
<GID>56</GID>
<name>OUT_6</name></connection>
<intersection>-117 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-33,-117,-6,-117</points>
<intersection>-33 0</intersection>
<intersection>-6 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-6,-118.5,-6,-117</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>-117 3</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,-106,-52,-106</points>
<connection>
<GID>85</GID>
<name>N_in0</name></connection>
<intersection>-71 6</intersection>
<intersection>-68 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-68,-111.5,-68,-106</points>
<intersection>-111.5 5</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-68,-111.5,-56,-111.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-68 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-71,-156,-71,-106</points>
<intersection>-156 8</intersection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>177,-156,177,49.5</points>
<intersection>-156 8</intersection>
<intersection>5 34</intersection>
<intersection>49.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-73.5,-156,177,-156</points>
<connection>
<GID>30</GID>
<name>N_in1</name></connection>
<intersection>-71 6</intersection>
<intersection>-41.5 13</intersection>
<intersection>-34 11</intersection>
<intersection>-19.5 31</intersection>
<intersection>4.5 12</intersection>
<intersection>123.5 29</intersection>
<intersection>177 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-106.5,49.5,177,49.5</points>
<connection>
<GID>28</GID>
<name>N_in1</name></connection>
<intersection>-87.5 15</intersection>
<intersection>-22 10</intersection>
<intersection>64 21</intersection>
<intersection>177 7</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-22,-10,-22,49.5</points>
<connection>
<GID>62</GID>
<name>OUT_7</name></connection>
<intersection>49.5 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-34,-156,-34,-148</points>
<connection>
<GID>56</GID>
<name>IN_7</name></connection>
<intersection>-156 8</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>4.5,-161,4.5,-156</points>
<connection>
<GID>2</GID>
<name>IN_7</name></connection>
<intersection>-156 8</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-41.5,-157,-41.5,-156</points>
<connection>
<GID>22</GID>
<name>OUT_7</name></connection>
<intersection>-156 8</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-87.5,-13,-87.5,49.5</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>49.5 9</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>64,4.5,64,49.5</points>
<intersection>4.5 24</intersection>
<intersection>49.5 9</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>91.5,-25.5,91.5,19.5</points>
<connection>
<GID>232</GID>
<name>IN_7</name></connection>
<connection>
<GID>231</GID>
<name>IN_7</name></connection>
<connection>
<GID>230</GID>
<name>IN_7</name></connection>
<connection>
<GID>229</GID>
<name>IN_7</name></connection>
<intersection>4.5 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>64,4.5,91.5,4.5</points>
<intersection>64 21</intersection>
<intersection>91.5 22</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>123.5,-156,123.5,-115</points>
<connection>
<GID>333</GID>
<name>N_in2</name></connection>
<intersection>-156 8</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-19.5,-182,-19.5,-156</points>
<intersection>-182 35</intersection>
<intersection>-156 8</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>169.5,5,177,5</points>
<connection>
<GID>225</GID>
<name>OUT_7</name></connection>
<intersection>177 7</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>-19.5,-182,-18,-182</points>
<connection>
<GID>73</GID>
<name>IN_7</name></connection>
<intersection>-19.5 31</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-111.5,-52,-111.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-112.5,-52,-112.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-114.5,-52,-114.5</points>
<connection>
<GID>83</GID>
<name>IN_3</name></connection>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-113.5,-52,-113.5</points>
<connection>
<GID>83</GID>
<name>IN_2</name></connection>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-115.5,-52,-115.5</points>
<connection>
<GID>83</GID>
<name>IN_4</name></connection>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-116.5,-52,-116.5</points>
<connection>
<GID>83</GID>
<name>IN_5</name></connection>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-117.5,-52,-117.5</points>
<connection>
<GID>83</GID>
<name>IN_6</name></connection>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-118.5,-52,-118.5</points>
<connection>
<GID>83</GID>
<name>IN_7</name></connection>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-114,-57,-112.5</points>
<intersection>-114 1</intersection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,-114,-57,-114</points>
<intersection>-71 3</intersection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-112.5,-56,-112.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-71,-155,-71,-114</points>
<intersection>-155 7</intersection>
<intersection>-114 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>176,-155,176,48.5</points>
<intersection>-155 7</intersection>
<intersection>4 35</intersection>
<intersection>48.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-155,176,-155</points>
<connection>
<GID>34</GID>
<name>N_in1</name></connection>
<intersection>-71 3</intersection>
<intersection>-40.5 15</intersection>
<intersection>-33 12</intersection>
<intersection>-20 33</intersection>
<intersection>3.5 13</intersection>
<intersection>126.5 30</intersection>
<intersection>176 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,48.5,176,48.5</points>
<connection>
<GID>33</GID>
<name>N_in1</name></connection>
<intersection>-88.5 16</intersection>
<intersection>-21 9</intersection>
<intersection>65.5 22</intersection>
<intersection>176 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-21,-10,-21,48.5</points>
<connection>
<GID>62</GID>
<name>OUT_6</name></connection>
<intersection>48.5 8</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-33,-155,-33,-148</points>
<connection>
<GID>56</GID>
<name>IN_6</name></connection>
<intersection>-155 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>3.5,-161,3.5,-155</points>
<connection>
<GID>2</GID>
<name>IN_6</name></connection>
<intersection>-155 7</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-40.5,-157,-40.5,-155</points>
<connection>
<GID>22</GID>
<name>OUT_6</name></connection>
<intersection>-155 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-88.5,-13,-88.5,48.5</points>
<connection>
<GID>209</GID>
<name>OUT_1</name></connection>
<intersection>48.5 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>65.5,1.5,65.5,48.5</points>
<intersection>1.5 25</intersection>
<intersection>48.5 8</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>91.5,-26.5,91.5,18.5</points>
<connection>
<GID>232</GID>
<name>IN_6</name></connection>
<connection>
<GID>231</GID>
<name>IN_6</name></connection>
<connection>
<GID>230</GID>
<name>IN_6</name></connection>
<connection>
<GID>229</GID>
<name>IN_6</name></connection>
<intersection>1.5 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>65.5,1.5,91.5,1.5</points>
<intersection>65.5 22</intersection>
<intersection>91.5 23</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>126.5,-155,126.5,-115</points>
<connection>
<GID>334</GID>
<name>N_in2</name></connection>
<intersection>-155 7</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>-20,-183,-20,-155</points>
<intersection>-183 36</intersection>
<intersection>-155 7</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>169.5,4,176,4</points>
<connection>
<GID>225</GID>
<name>OUT_6</name></connection>
<intersection>176 6</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>-20,-183,-18,-183</points>
<connection>
<GID>73</GID>
<name>IN_6</name></connection>
<intersection>-20 33</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-113.5,-57,-111.5</points>
<intersection>-113.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,-111.5,-57,-111.5</points>
<intersection>-68.5 3</intersection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-113.5,-56,-113.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-68.5,-112,-68.5,-111.5</points>
<intersection>-112 4</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-71,-112,-68.5,-112</points>
<intersection>-71 5</intersection>
<intersection>-68.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-71,-154,-71,-112</points>
<intersection>-154 7</intersection>
<intersection>-112 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>175,-154,175,47.5</points>
<intersection>-154 7</intersection>
<intersection>3 33</intersection>
<intersection>47.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-154,175,-154</points>
<connection>
<GID>36</GID>
<name>N_in1</name></connection>
<intersection>-71 5</intersection>
<intersection>-39.5 13</intersection>
<intersection>-32 10</intersection>
<intersection>-20.5 31</intersection>
<intersection>2.5 11</intersection>
<intersection>129.5 28</intersection>
<intersection>175 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,47.5,175,47.5</points>
<connection>
<GID>35</GID>
<name>N_in1</name></connection>
<intersection>-89.5 14</intersection>
<intersection>-20 9</intersection>
<intersection>67 20</intersection>
<intersection>175 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-20,-10,-20,47.5</points>
<connection>
<GID>62</GID>
<name>OUT_5</name></connection>
<intersection>47.5 8</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-32,-154,-32,-148</points>
<connection>
<GID>56</GID>
<name>IN_5</name></connection>
<intersection>-154 7</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>2.5,-161,2.5,-154</points>
<connection>
<GID>2</GID>
<name>IN_5</name></connection>
<intersection>-154 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-39.5,-157,-39.5,-154</points>
<connection>
<GID>22</GID>
<name>OUT_5</name></connection>
<intersection>-154 7</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-89.5,-13,-89.5,47.5</points>
<connection>
<GID>209</GID>
<name>OUT_2</name></connection>
<intersection>47.5 8</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>67,-1.5,67,47.5</points>
<intersection>-1.5 23</intersection>
<intersection>47.5 8</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>91.5,-27.5,91.5,17.5</points>
<connection>
<GID>232</GID>
<name>IN_5</name></connection>
<connection>
<GID>231</GID>
<name>IN_5</name></connection>
<connection>
<GID>230</GID>
<name>IN_5</name></connection>
<connection>
<GID>229</GID>
<name>IN_5</name></connection>
<intersection>-1.5 23</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>67,-1.5,91.5,-1.5</points>
<intersection>67 20</intersection>
<intersection>91.5 21</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>129.5,-154,129.5,-115</points>
<connection>
<GID>335</GID>
<name>N_in2</name></connection>
<intersection>-154 7</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-20.5,-184,-20.5,-154</points>
<intersection>-184 34</intersection>
<intersection>-154 7</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>169.5,3,175,3</points>
<connection>
<GID>225</GID>
<name>OUT_5</name></connection>
<intersection>175 6</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>-20.5,-184,-18,-184</points>
<connection>
<GID>73</GID>
<name>IN_5</name></connection>
<intersection>-20.5 31</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-114.5,-57,-111.5</points>
<intersection>-114.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-111.5,-57,-111.5</points>
<intersection>-68 3</intersection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-114.5,-56,-114.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-68,-115,-68,-111.5</points>
<intersection>-115 4</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-71,-115,-68,-115</points>
<intersection>-71 5</intersection>
<intersection>-68 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-71,-153,-71,-115</points>
<intersection>-153 7</intersection>
<intersection>-115 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>174,-153,174,46.5</points>
<intersection>-153 7</intersection>
<intersection>2 36</intersection>
<intersection>46.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-153,174,-153</points>
<connection>
<GID>38</GID>
<name>N_in1</name></connection>
<intersection>-71 5</intersection>
<intersection>-38.5 14</intersection>
<intersection>-31 11</intersection>
<intersection>1.5 12</intersection>
<intersection>132.5 29</intersection>
<intersection>174 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,46.5,174,46.5</points>
<connection>
<GID>37</GID>
<name>N_in1</name></connection>
<intersection>-90.5 15</intersection>
<intersection>-19 9</intersection>
<intersection>68.5 21</intersection>
<intersection>174 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-19,-10,-19,46.5</points>
<connection>
<GID>62</GID>
<name>OUT_4</name></connection>
<intersection>46.5 8</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-31,-153,-31,-148</points>
<connection>
<GID>56</GID>
<name>IN_4</name></connection>
<intersection>-153 7</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>1.5,-179.5,1.5,-153</points>
<connection>
<GID>2</GID>
<name>IN_4</name></connection>
<intersection>-179.5 33</intersection>
<intersection>-153 7</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-38.5,-157,-38.5,-153</points>
<connection>
<GID>22</GID>
<name>OUT_4</name></connection>
<intersection>-153 7</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-90.5,-13,-90.5,46.5</points>
<connection>
<GID>209</GID>
<name>OUT_3</name></connection>
<intersection>46.5 8</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>68.5,-4.5,68.5,46.5</points>
<intersection>-4.5 24</intersection>
<intersection>46.5 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>91.5,-28.5,91.5,16.5</points>
<connection>
<GID>232</GID>
<name>IN_4</name></connection>
<connection>
<GID>231</GID>
<name>IN_4</name></connection>
<connection>
<GID>230</GID>
<name>IN_4</name></connection>
<connection>
<GID>229</GID>
<name>IN_4</name></connection>
<intersection>-4.5 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>68.5,-4.5,91.5,-4.5</points>
<intersection>68.5 21</intersection>
<intersection>91.5 22</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>132.5,-153,132.5,-115</points>
<connection>
<GID>336</GID>
<name>N_in2</name></connection>
<intersection>-153 7</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-18,-179.5,1.5,-179.5</points>
<intersection>-18 34</intersection>
<intersection>1.5 12</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>-18,-185,-18,-179.5</points>
<connection>
<GID>73</GID>
<name>IN_4</name></connection>
<intersection>-179.5 33</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>169.5,2,174,2</points>
<connection>
<GID>225</GID>
<name>OUT_4</name></connection>
<intersection>174 6</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-115.5,-57,-111.5</points>
<intersection>-115.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,-111.5,-57,-111.5</points>
<intersection>-68 3</intersection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-115.5,-56,-115.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-68,-118,-68,-111.5</points>
<intersection>-118 4</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-69.5,-118,-68,-118</points>
<intersection>-69.5 5</intersection>
<intersection>-68 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-69.5,-152,-69.5,-118</points>
<intersection>-152 7</intersection>
<intersection>-118 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>173,-152,173,45.5</points>
<intersection>-152 7</intersection>
<intersection>1 38</intersection>
<intersection>45.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-152,173,-152</points>
<connection>
<GID>40</GID>
<name>N_in1</name></connection>
<intersection>-69.5 5</intersection>
<intersection>-37.5 15</intersection>
<intersection>-30 12</intersection>
<intersection>-21.5 13</intersection>
<intersection>135.5 32</intersection>
<intersection>173 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,45.5,173,45.5</points>
<connection>
<GID>39</GID>
<name>N_in1</name></connection>
<intersection>-91.5 16</intersection>
<intersection>-18 10</intersection>
<intersection>69.5 24</intersection>
<intersection>173 6</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-18,-10,-18,45.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>45.5 8</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-30,-152,-30,-148</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>-152 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-21.5,-180,-21.5,-152</points>
<intersection>-180 35</intersection>
<intersection>-161 39</intersection>
<intersection>-152 7</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-37.5,-157,-37.5,-152</points>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<intersection>-152 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-91.5,-13,-91.5,45.5</points>
<connection>
<GID>209</GID>
<name>OUT_4</name></connection>
<intersection>45.5 8</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>69.5,-7.5,69.5,45.5</points>
<intersection>-7.5 27</intersection>
<intersection>45.5 8</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>91.5,-29.5,91.5,15.5</points>
<connection>
<GID>232</GID>
<name>IN_3</name></connection>
<connection>
<GID>231</GID>
<name>IN_3</name></connection>
<connection>
<GID>230</GID>
<name>IN_3</name></connection>
<connection>
<GID>229</GID>
<name>IN_3</name></connection>
<intersection>-7.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>69.5,-7.5,91.5,-7.5</points>
<intersection>69.5 24</intersection>
<intersection>91.5 25</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>135.5,-152,135.5,-115</points>
<connection>
<GID>337</GID>
<name>N_in2</name></connection>
<intersection>-152 7</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>-21.5,-180,-18,-180</points>
<intersection>-21.5 13</intersection>
<intersection>-18 36</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>-18,-186,-18,-180</points>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<intersection>-180 35</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>169.5,1,173,1</points>
<connection>
<GID>225</GID>
<name>OUT_3</name></connection>
<intersection>173 6</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-21.5,-161,0.5,-161</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>-21.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-116.5,-57,-111.5</points>
<intersection>-116.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-111.5,-57,-111.5</points>
<intersection>-67.5 3</intersection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-116.5,-56,-116.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-67.5,-121,-67.5,-111.5</points>
<intersection>-121 4</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-70,-121,-67.5,-121</points>
<intersection>-70 5</intersection>
<intersection>-67.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-70,-151,-70,-121</points>
<intersection>-151 7</intersection>
<intersection>-121 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>172,-151,172,44.5</points>
<intersection>-151 7</intersection>
<intersection>0 38</intersection>
<intersection>44.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-151,172,-151</points>
<connection>
<GID>42</GID>
<name>N_in1</name></connection>
<intersection>-70 5</intersection>
<intersection>-36.5 16</intersection>
<intersection>-29 13</intersection>
<intersection>-17 14</intersection>
<intersection>138.5 32</intersection>
<intersection>172 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,44.5,172,44.5</points>
<connection>
<GID>41</GID>
<name>N_in1</name></connection>
<intersection>-92.5 17</intersection>
<intersection>-17 12</intersection>
<intersection>70 22</intersection>
<intersection>172 6</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-17,-10,-17,44.5</points>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection>
<intersection>44.5 8</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-29,-151,-29,-148</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>-151 7</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-17,-187,-17,-151</points>
<intersection>-187 40</intersection>
<intersection>-161 39</intersection>
<intersection>-151 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-36.5,-157,-36.5,-151</points>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<intersection>-151 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-92.5,-13,-92.5,44.5</points>
<connection>
<GID>209</GID>
<name>OUT_5</name></connection>
<intersection>44.5 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>70,-10.5,70,44.5</points>
<intersection>-10.5 25</intersection>
<intersection>44.5 8</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>91.5,-30.5,91.5,14.5</points>
<connection>
<GID>232</GID>
<name>IN_2</name></connection>
<connection>
<GID>231</GID>
<name>IN_2</name></connection>
<connection>
<GID>230</GID>
<name>IN_2</name></connection>
<connection>
<GID>229</GID>
<name>IN_2</name></connection>
<intersection>-10.5 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>70,-10.5,91.5,-10.5</points>
<intersection>70 22</intersection>
<intersection>91.5 23</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>138.5,-151,138.5,-115</points>
<connection>
<GID>338</GID>
<name>N_in2</name></connection>
<intersection>-151 7</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>169.5,0,172,0</points>
<connection>
<GID>225</GID>
<name>OUT_2</name></connection>
<intersection>172 6</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-17,-161,-0.5,-161</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-17 14</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>-18,-187,-17,-187</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>-17 14</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-117.5,-57,-111.5</points>
<intersection>-117.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,-111.5,-57,-111.5</points>
<intersection>-66.5 3</intersection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-117.5,-56,-117.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-66.5,-124,-66.5,-111.5</points>
<intersection>-124 4</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-70.5,-124,-66.5,-124</points>
<intersection>-70.5 5</intersection>
<intersection>-66.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-70.5,-150,-70.5,-124</points>
<intersection>-150 7</intersection>
<intersection>-124 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>171,-150,171,43.5</points>
<intersection>-150 7</intersection>
<intersection>-1 36</intersection>
<intersection>43.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-150,171,-150</points>
<connection>
<GID>44</GID>
<name>N_in1</name></connection>
<intersection>-70.5 5</intersection>
<intersection>-35.5 15</intersection>
<intersection>-28 11</intersection>
<intersection>-14 12</intersection>
<intersection>141.5 30</intersection>
<intersection>171 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,43.5,171,43.5</points>
<connection>
<GID>43</GID>
<name>N_in1</name></connection>
<intersection>-93.5 16</intersection>
<intersection>-16 10</intersection>
<intersection>71.5 21</intersection>
<intersection>171 6</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-16,-10,-16,43.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<intersection>43.5 8</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-28,-150,-28,-148</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-150 7</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-14,-172,-14,-150</points>
<intersection>-172 33</intersection>
<intersection>-161 38</intersection>
<intersection>-150 7</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-35.5,-157,-35.5,-150</points>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<intersection>-150 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-93.5,-13,-93.5,43.5</points>
<connection>
<GID>209</GID>
<name>OUT_6</name></connection>
<intersection>43.5 8</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>71.5,-13.5,71.5,43.5</points>
<intersection>-13.5 24</intersection>
<intersection>43.5 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>91.5,-31.5,91.5,13.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>-13.5 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>71.5,-13.5,91.5,-13.5</points>
<intersection>71.5 21</intersection>
<intersection>91.5 22</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>141.5,-150,141.5,-115</points>
<connection>
<GID>339</GID>
<name>N_in2</name></connection>
<intersection>-150 7</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-19,-172,-14,-172</points>
<intersection>-19 34</intersection>
<intersection>-14 12</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>-19,-188,-19,-172</points>
<intersection>-188 37</intersection>
<intersection>-172 33</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>169.5,-1,171,-1</points>
<connection>
<GID>225</GID>
<name>OUT_1</name></connection>
<intersection>171 6</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-19,-188,-18,-188</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>-19 34</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>-14,-161,-1.5,-161</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-14 12</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-118.5,-57,-111.5</points>
<intersection>-118.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,-111.5,-57,-111.5</points>
<intersection>-65.5 3</intersection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-118.5,-56,-118.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-65.5,-127,-65.5,-111.5</points>
<intersection>-127 4</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-71,-127,-65.5,-127</points>
<intersection>-71 5</intersection>
<intersection>-65.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-71,-149,-71,-127</points>
<intersection>-149 7</intersection>
<intersection>-127 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>170,-149,170,42.5</points>
<intersection>-149 7</intersection>
<intersection>-2 38</intersection>
<intersection>42.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-73.5,-149,170,-149</points>
<connection>
<GID>46</GID>
<name>N_in1</name></connection>
<intersection>-71 5</intersection>
<intersection>-34.5 16</intersection>
<intersection>-27 12</intersection>
<intersection>-13.5 13</intersection>
<intersection>144.5 31</intersection>
<intersection>170 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,42.5,170,42.5</points>
<connection>
<GID>45</GID>
<name>N_in1</name></connection>
<intersection>-94.5 17</intersection>
<intersection>-15 11</intersection>
<intersection>72.5 22</intersection>
<intersection>170 6</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-15,-10,-15,42.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>42.5 8</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-27,-149,-27,-148</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-149 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-13.5,-172.5,-13.5,-149</points>
<intersection>-172.5 34</intersection>
<intersection>-161 39</intersection>
<intersection>-149 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-34.5,-157,-34.5,-149</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-149 7</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-94.5,-13,-94.5,42.5</points>
<connection>
<GID>209</GID>
<name>OUT_7</name></connection>
<intersection>42.5 8</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>72.5,-16.5,72.5,42.5</points>
<intersection>-16.5 25</intersection>
<intersection>42.5 8</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>91.5,-32.5,91.5,12.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>-16.5 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>72.5,-16.5,91.5,-16.5</points>
<intersection>72.5 22</intersection>
<intersection>91.5 23</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>144.5,-149,144.5,-115</points>
<connection>
<GID>340</GID>
<name>N_in2</name></connection>
<intersection>-149 7</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>-18.5,-172.5,-13.5,-172.5</points>
<intersection>-18.5 35</intersection>
<intersection>-13.5 13</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>-18.5,-189,-18.5,-172.5</points>
<intersection>-189 40</intersection>
<intersection>-172.5 34</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>169.5,-2,170,-2</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>170 6</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>-13.5,-161,-2.5,-161</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-13.5 13</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>-18.5,-189,-18,-189</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-18.5 35</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-115,-46,-115</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<connection>
<GID>95</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-111.5,-33,-111.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-115,-42.5,-79</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-115 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42.5,-111.5,-37,-111.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44,-115,-42.5,-115</points>
<connection>
<GID>95</GID>
<name>N_in1</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43.5,-109.5,-43.5,-106</points>
<intersection>-109.5 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43.5,-109.5,-37,-109.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-58,-106,-43.5,-106</points>
<connection>
<GID>85</GID>
<name>N_in1</name></connection>
<intersection>-58 4</intersection>
<intersection>-43.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-58,-106,-58,-79</points>
<intersection>-106 2</intersection>
<intersection>-79 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-58,-79,-57.5,-79</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-58 4</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-34.5,-105,-23,-105</points>
<connection>
<GID>100</GID>
<name>N_in0</name></connection>
<intersection>-34.5 4</intersection>
<intersection>-27 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-34.5,-105,-34.5,-79</points>
<intersection>-105 1</intersection>
<intersection>-79 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-27,-110.5,-27,-105</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-34.5,-79,-29,-79</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-34.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-109.5,-33,-109.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-79,-23,-75.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,-75.5,-23,-75.5</points>
<connection>
<GID>110</GID>
<name>N_in1</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-79,-36.5,-75.5</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-38,-75.5,-36.5,-75.5</points>
<connection>
<GID>109</GID>
<name>N_in1</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,-90.5,-30,-90.5</points>
<intersection>-58 15</intersection>
<intersection>-42.5 16</intersection>
<intersection>-30 17</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-58,-90.5,-58,-81.5</points>
<intersection>-90.5 1</intersection>
<intersection>-81.5 19</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-42.5,-90.5,-42.5,-83</points>
<connection>
<GID>112</GID>
<name>clock_enable</name></connection>
<intersection>-90.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-30,-90.5,-30,-81.5</points>
<intersection>-90.5 1</intersection>
<intersection>-81.5 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-58,-81.5,38,-81.5</points>
<intersection>-58 15</intersection>
<intersection>-57.5 24</intersection>
<intersection>-30 17</intersection>
<intersection>-29 25</intersection>
<intersection>38 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>38,-143.5,38,-81.5</points>
<intersection>-143.5 26</intersection>
<intersection>-81.5 19</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>-57.5,-83,-57.5,-81.5</points>
<connection>
<GID>102</GID>
<name>clock_enable</name></connection>
<intersection>-81.5 19</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>-29,-83,-29,-81.5</points>
<connection>
<GID>114</GID>
<name>clock_enable</name></connection>
<intersection>-81.5 19</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>30.5,-143.5,38,-143.5</points>
<intersection>30.5 27</intersection>
<intersection>38 23</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>30.5,-143.5,30.5,-142</points>
<intersection>-143.5 26</intersection>
<intersection>-142 29</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>30,-142,30.5,-142</points>
<connection>
<GID>135</GID>
<name>OUT_1</name></connection>
<intersection>30.5 27</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-79,-51.5,-75.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-52,-75.5,-51.5,-75.5</points>
<connection>
<GID>108</GID>
<name>N_in1</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40.5,-71.5,-40.5,-68.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-39,-74.5,-39,-71.5</points>
<connection>
<GID>109</GID>
<name>N_in3</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-40.5,-71.5,-39,-71.5</points>
<intersection>-40.5 0</intersection>
<intersection>-39 1</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,-71.5,-54,-68.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-53,-74.5,-53,-71.5</points>
<connection>
<GID>108</GID>
<name>N_in3</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-54,-71.5,-53,-71.5</points>
<intersection>-54 0</intersection>
<intersection>-53 1</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-71.5,-27,-68.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-25.5,-74.5,-25.5,-71.5</points>
<connection>
<GID>110</GID>
<name>N_in3</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-27,-71.5,-25.5,-71.5</points>
<intersection>-27 0</intersection>
<intersection>-25.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-72.5,4.5,-62.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-26,-62.5,4.5,-62.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-72.5,2.5,-61.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-39.5,-61.5,2.5,-61.5</points>
<intersection>-39.5 3</intersection>
<intersection>2.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-39.5,-62.5,-39.5,-61.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-61.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>0.5,-72.5,0.5,-60.5</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-53,-60.5,0.5,-60.5</points>
<intersection>-53 3</intersection>
<intersection>0.5 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-53,-62.5,-53,-60.5</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>-60.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-104,-46.5,22.5</points>
<intersection>-104 2</intersection>
<intersection>-68.5 3</intersection>
<intersection>22.5 10</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-40,-138.5,-40,-96</points>
<intersection>-138.5 4</intersection>
<intersection>-104 2</intersection>
<intersection>-96 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-46.5,-104,-40,-104</points>
<intersection>-46.5 0</intersection>
<intersection>-40 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-52,-68.5,-46.5,-68.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-46.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-40,-138.5,-32,-138.5</points>
<intersection>-40 1</intersection>
<intersection>-32 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-32,-140,-32,-138.5</points>
<connection>
<GID>56</GID>
<name>OUT_5</name></connection>
<intersection>-138.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-40,-96,-14.5,-96</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>-40 1</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-46.5,22.5,45,22.5</points>
<intersection>-46.5 0</intersection>
<intersection>45 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>45,22.5,45,31.5</points>
<intersection>22.5 10</intersection>
<intersection>31.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>45,31.5,80,31.5</points>
<connection>
<GID>226</GID>
<name>N_in0</name></connection>
<intersection>45 11</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-99.5,-35.5,27.5</points>
<intersection>-99.5 2</intersection>
<intersection>-68.5 3</intersection>
<intersection>27.5 5</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-31,-140,-31,-99.5</points>
<connection>
<GID>56</GID>
<name>OUT_4</name></connection>
<intersection>-99.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-35.5,-99.5,-31,-99.5</points>
<intersection>-35.5 0</intersection>
<intersection>-31 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-38.5,-68.5,-35.5,-68.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-35.5,27.5,100,27.5</points>
<connection>
<GID>227</GID>
<name>N_in0</name></connection>
<intersection>-35.5 0</intersection>
<intersection>100 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>100,27.5,100,28</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>27.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21.5,-102.5,-21.5,-68.5</points>
<intersection>-102.5 2</intersection>
<intersection>-68.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-30,-140,-30,30.5</points>
<connection>
<GID>56</GID>
<name>OUT_3</name></connection>
<intersection>-102.5 2</intersection>
<intersection>-54 4</intersection>
<intersection>30.5 14</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,-102.5,-21.5,-102.5</points>
<intersection>-30 1</intersection>
<intersection>-21.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-25,-68.5,-21.5,-68.5</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-21.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-98,-54,-30,-54</points>
<intersection>-98 9</intersection>
<intersection>-95 10</intersection>
<intersection>-92 11</intersection>
<intersection>-89 12</intersection>
<intersection>-86 13</intersection>
<intersection>-30 1</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-98,-54,-98,-50.5</points>
<connection>
<GID>153</GID>
<name>N_in2</name></connection>
<intersection>-54 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-95,-54,-95,-50.5</points>
<connection>
<GID>154</GID>
<name>N_in2</name></connection>
<intersection>-54 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-92,-54,-92,-50.5</points>
<connection>
<GID>155</GID>
<name>N_in2</name></connection>
<intersection>-54 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-89,-54,-89,-50.5</points>
<connection>
<GID>156</GID>
<name>N_in2</name></connection>
<intersection>-54 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-86,-54,-86,-50.5</points>
<connection>
<GID>157</GID>
<name>N_in2</name></connection>
<intersection>-54 4</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-30,30.5,100,30.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>-30 1</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-27,-140,-27,26.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 2</intersection>
<intersection>26.5 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-77,-59.5,-27,-59.5</points>
<intersection>-77 7</intersection>
<intersection>-59 3</intersection>
<intersection>-27 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-59,-59.5,-59,-56</points>
<connection>
<GID>150</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-77,-59.5,-77,-50.5</points>
<connection>
<GID>160</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-27,26.5,113.5,26.5</points>
<intersection>-27 1</intersection>
<intersection>113.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>113.5,26.5,113.5,28.5</points>
<intersection>26.5 8</intersection>
<intersection>28.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>113,28.5,113.5,28.5</points>
<connection>
<GID>281</GID>
<name>N_in1</name></connection>
<intersection>113.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-59.5,-62,-56</points>
<connection>
<GID>149</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-28,-140,-28,36</points>
<connection>
<GID>56</GID>
<name>OUT_1</name></connection>
<intersection>-59.5 2</intersection>
<intersection>36 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-80,-59.5,-28,-59.5</points>
<intersection>-80 4</intersection>
<intersection>-62 0</intersection>
<intersection>-28 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-80,-59.5,-80,-50.5</points>
<connection>
<GID>159</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-28,36,114,36</points>
<intersection>-28 1</intersection>
<intersection>114 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>114,31.5,114,36</points>
<intersection>31.5 9</intersection>
<intersection>36 5</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>113,31.5,114,31.5</points>
<connection>
<GID>279</GID>
<name>N_in1</name></connection>
<intersection>114 8</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-59.5,-65,-56</points>
<connection>
<GID>148</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-29,-140,-29,26</points>
<connection>
<GID>56</GID>
<name>OUT_2</name></connection>
<intersection>-59.5 2</intersection>
<intersection>26 15</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-83,-59.5,-29,-59.5</points>
<intersection>-83 14</intersection>
<intersection>-81 8</intersection>
<intersection>-77.5 9</intersection>
<intersection>-74 10</intersection>
<intersection>-71 11</intersection>
<intersection>-68 12</intersection>
<intersection>-65 0</intersection>
<intersection>-29 1</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-81,-59.5,-81,-56</points>
<connection>
<GID>142</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-77.5,-59.5,-77.5,-56</points>
<connection>
<GID>143</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-74,-59.5,-74,-56</points>
<connection>
<GID>145</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-71,-59.5,-71,-56</points>
<connection>
<GID>146</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-68,-59.5,-68,-56</points>
<connection>
<GID>147</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-83,-59.5,-83,-50.5</points>
<connection>
<GID>158</GID>
<name>N_in2</name></connection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-29,26,100,26</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>29,-75.5,32,-75.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-75.5,32,-74</points>
<connection>
<GID>127</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-75.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>30,-74,31,-74</points>
<connection>
<GID>127</GID>
<name>DATA_OUT_1</name></connection>
<intersection>30 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>30,-75.5,30,-74</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>-74 7</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30,-75.5,31,-75.5</points>
<connection>
<GID>121</GID>
<name>IN_2</name></connection>
<intersection>30 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-75.5,30,-74</points>
<connection>
<GID>127</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-75.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>29,-75.5,32,-75.5</points>
<connection>
<GID>121</GID>
<name>IN_3</name></connection>
<intersection>29 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29,-75.5,29,-74</points>
<connection>
<GID>127</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-75.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-38.5,51.5,-38.5</points>
<intersection>-106 72</intersection>
<intersection>-101 71</intersection>
<intersection>-96 70</intersection>
<intersection>-91 69</intersection>
<intersection>-86 68</intersection>
<intersection>-81 67</intersection>
<intersection>-76 66</intersection>
<intersection>-71 65</intersection>
<intersection>51.5 58</intersection></hsegment>
<vsegment>
<ID>58</ID>
<points>51.5,-126.5,51.5,-38.5</points>
<intersection>-126.5 61</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>61</ID>
<points>51.5,-126.5,55.5,-126.5</points>
<intersection>51.5 58</intersection>
<intersection>55.5 62</intersection></hsegment>
<vsegment>
<ID>62</ID>
<points>55.5,-126.5,55.5,-122.5</points>
<intersection>-126.5 61</intersection>
<intersection>-122.5 63</intersection></vsegment>
<hsegment>
<ID>63</ID>
<points>55.5,-122.5,56,-122.5</points>
<intersection>55.5 62</intersection>
<intersection>56 64</intersection></hsegment>
<vsegment>
<ID>64</ID>
<points>56,-124,56,-122.5</points>
<connection>
<GID>140</GID>
<name>OUT_3</name></connection>
<intersection>-122.5 63</intersection></vsegment>
<vsegment>
<ID>65</ID>
<points>-71,-41,-71,-38.5</points>
<connection>
<GID>172</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>66</ID>
<points>-76,-41,-76,-38.5</points>
<connection>
<GID>171</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>67</ID>
<points>-81,-41,-81,-38.5</points>
<connection>
<GID>170</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>68</ID>
<points>-86,-41,-86,-38.5</points>
<connection>
<GID>169</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>69</ID>
<points>-91,-41,-91,-38.5</points>
<connection>
<GID>168</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>70</ID>
<points>-96,-41,-96,-38.5</points>
<connection>
<GID>167</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>71</ID>
<points>-101,-41,-101,-38.5</points>
<connection>
<GID>166</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>72</ID>
<points>-106,-41,-106,-38.5</points>
<connection>
<GID>165</GID>
<name>SEL_0</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-78.5,35,-78.5</points>
<connection>
<GID>121</GID>
<name>load</name></connection>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-94,32,-93.5</points>
<connection>
<GID>129</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-94 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,-94.5,29,-94</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29,-94,32,-94</points>
<intersection>29 1</intersection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-94,31,-93.5</points>
<connection>
<GID>129</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-94 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30,-94.5,30,-94</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30,-94,31,-94</points>
<intersection>30 1</intersection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-94,30,-93.5</points>
<connection>
<GID>129</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-94 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,-94.5,31,-94</points>
<connection>
<GID>124</GID>
<name>IN_2</name></connection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30,-94,31,-94</points>
<intersection>30 0</intersection>
<intersection>31 1</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-86.5,-32.5,-84,-32.5</points>
<connection>
<GID>174</GID>
<name>carry_out</name></connection>
<connection>
<GID>175</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-94,29,-93.5</points>
<connection>
<GID>129</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-94 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32,-94.5,32,-94</points>
<connection>
<GID>124</GID>
<name>IN_3</name></connection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29,-94,32,-94</points>
<intersection>29 0</intersection>
<intersection>32 1</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>35.5,-69.5,35.5,-69.5</points>
<connection>
<GID>127</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-89,35.5,-89</points>
<connection>
<GID>129</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>274</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>35,-109,35,-109</points>
<connection>
<GID>131</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-128.5,35.5,-128.5</points>
<connection>
<GID>276</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-88.5,59.5,-88.5</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<connection>
<GID>295</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-54,-67.5,-43</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-67.5,-54,-59,-54</points>
<connection>
<GID>150</GID>
<name>N_in3</name></connection>
<intersection>-67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,-54,-72.5,-43</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-72.5,-54,-62,-54</points>
<connection>
<GID>149</GID>
<name>N_in3</name></connection>
<intersection>-72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-77.5,-54,-77.5,-43</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-54,-65,-54</points>
<connection>
<GID>148</GID>
<name>N_in3</name></connection>
<intersection>-77.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82.5,-54,-82.5,-43</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-82.5,-54,-68,-54</points>
<connection>
<GID>147</GID>
<name>N_in3</name></connection>
<intersection>-82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-87.5,-54,-87.5,-43</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-54,-71,-54</points>
<connection>
<GID>146</GID>
<name>N_in3</name></connection>
<intersection>-87.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92.5,-54,-92.5,-43</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-92.5,-54,-74,-54</points>
<connection>
<GID>145</GID>
<name>N_in3</name></connection>
<intersection>-92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-97.5,-54,-97.5,-43</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-97.5,-54,-77.5,-54</points>
<connection>
<GID>143</GID>
<name>N_in3</name></connection>
<intersection>-97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-102.5,-54,-102.5,-43</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-102.5,-54,-81,-54</points>
<connection>
<GID>142</GID>
<name>N_in3</name></connection>
<intersection>-102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-51.5,-69.5,-43</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-77,-51.5,-77,-48.5</points>
<connection>
<GID>160</GID>
<name>N_in3</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-77,-51.5,-69.5,-51.5</points>
<intersection>-77 1</intersection>
<intersection>-69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,-52,-80,-48.5</points>
<connection>
<GID>159</GID>
<name>N_in3</name></connection>
<intersection>-52 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-74.5,-52,-74.5,-43</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-80,-52,-74.5,-52</points>
<intersection>-80 0</intersection>
<intersection>-74.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-79.5,-51.5,-79.5,-43</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-83,-51.5,-83,-48.5</points>
<connection>
<GID>158</GID>
<name>N_in3</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-83,-51.5,-79.5,-51.5</points>
<intersection>-83 1</intersection>
<intersection>-79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86,-51.5,-86,-48.5</points>
<connection>
<GID>157</GID>
<name>N_in3</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-84.5,-51.5,-84.5,-43</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-86,-51.5,-84.5,-51.5</points>
<intersection>-86 0</intersection>
<intersection>-84.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89.5,-51.5,-89.5,-43</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-89,-51.5,-89,-48.5</points>
<connection>
<GID>156</GID>
<name>N_in3</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-89.5,-51.5,-89,-51.5</points>
<intersection>-89.5 0</intersection>
<intersection>-89 1</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92,-51.5,-92,-48.5</points>
<connection>
<GID>155</GID>
<name>N_in3</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-94.5,-51.5,-94.5,-43</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-94.5,-51.5,-92,-51.5</points>
<intersection>-94.5 1</intersection>
<intersection>-92 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-95,-48.5,-95,-43</points>
<connection>
<GID>154</GID>
<name>N_in3</name></connection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-99.5,-43,-95,-43</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>-95 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-104.5,-51.5,-104.5,-43</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-98,-51.5,-98,-48.5</points>
<connection>
<GID>153</GID>
<name>N_in3</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-104.5,-51.5,-98,-51.5</points>
<intersection>-104.5 0</intersection>
<intersection>-98 1</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-99.5,-37,-99.5,-35.5</points>
<connection>
<GID>174</GID>
<name>IN_B_0</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-68.5,-39,-68.5,-37</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-99.5,-37,-68.5,-37</points>
<intersection>-99.5 0</intersection>
<intersection>-68.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73.5,-39,-73.5,-37</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-98.5,-37,-98.5,-35.5</points>
<connection>
<GID>174</GID>
<name>IN_B_1</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-98.5,-37,-73.5,-37</points>
<intersection>-98.5 1</intersection>
<intersection>-73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-97.5,-37,-97.5,-35.5</points>
<connection>
<GID>174</GID>
<name>IN_B_2</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-78.5,-39,-78.5,-37</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-97.5,-37,-78.5,-37</points>
<intersection>-97.5 0</intersection>
<intersection>-78.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96.5,-37,-96.5,-35.5</points>
<connection>
<GID>174</GID>
<name>IN_B_3</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-83.5,-39,-83.5,-37</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-96.5,-37,-83.5,-37</points>
<intersection>-96.5 0</intersection>
<intersection>-83.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,-37,-81,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_B_0</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-88.5,-39,-88.5,-37</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-88.5,-37,-81,-37</points>
<intersection>-88.5 1</intersection>
<intersection>-81 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,-37,-80,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_B_1</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-93.5,-39,-93.5,-37</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-93.5,-37,-80,-37</points>
<intersection>-93.5 1</intersection>
<intersection>-80 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-79,-37,-79,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_B_2</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-98.5,-39,-98.5,-37</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-98.5,-37,-79,-37</points>
<intersection>-98.5 1</intersection>
<intersection>-79 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-37,-78,-35.5</points>
<connection>
<GID>175</GID>
<name>IN_B_3</name></connection>
<intersection>-37 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-103.5,-39,-103.5,-37</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-103.5,-37,-78,-37</points>
<intersection>-103.5 1</intersection>
<intersection>-78 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-109,59.5,-109</points>
<connection>
<GID>278</GID>
<name>OUT_0</name></connection>
<connection>
<GID>296</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-97.5,35,-97.5</points>
<connection>
<GID>124</GID>
<name>load</name></connection>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-117,34.5,-117</points>
<connection>
<GID>132</GID>
<name>load</name></connection>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-114,28.5,-113.5</points>
<connection>
<GID>131</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-114,31.5,-114</points>
<connection>
<GID>132</GID>
<name>IN_3</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-114,31.5,-113.5</points>
<connection>
<GID>131</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-114,31.5,-114</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-114,30.5,-113.5</points>
<connection>
<GID>131</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-114,30.5,-114</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-114,29.5,-113.5</points>
<connection>
<GID>131</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-114,30.5,-114</points>
<connection>
<GID>132</GID>
<name>IN_2</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36,-43.5,55.5,-43.5</points>
<intersection>-36 20</intersection>
<intersection>-31 19</intersection>
<intersection>-26 18</intersection>
<intersection>-21 17</intersection>
<intersection>-16 16</intersection>
<intersection>-11 15</intersection>
<intersection>-6 22</intersection>
<intersection>-1 21</intersection>
<intersection>55.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>55.5,-120,55.5,-43.5</points>
<intersection>-120 13</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>54,-120,55.5,-120</points>
<intersection>54 14</intersection>
<intersection>55.5 10</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>54,-124,54,-120</points>
<connection>
<GID>140</GID>
<name>OUT_1</name></connection>
<intersection>-120 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-11,-43.5,-11,-41.5</points>
<connection>
<GID>192</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-16,-43.5,-16,-41.5</points>
<connection>
<GID>191</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-21,-43.5,-21,-41.5</points>
<connection>
<GID>190</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-26,-43.5,-26,-41.5</points>
<connection>
<GID>189</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-31,-43.5,-31,-41.5</points>
<connection>
<GID>188</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>-36,-43.5,-36,-41.5</points>
<connection>
<GID>187</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>-1,-43.5,-1,-41.5</points>
<connection>
<GID>194</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>-6,-43.5,-6,-41.5</points>
<connection>
<GID>193</GID>
<name>SEL_0</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-43.5,-34.5,-35.5</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-96,-35.5,-96,-17</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-17 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-96,-35.5,-34.5,-35.5</points>
<intersection>-96 1</intersection>
<intersection>-34.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-96,-17,-94.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_7</name></connection>
<intersection>-96 1</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-133.5,31.5,-133</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-133.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29,-134,29,-133.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29,-133.5,31.5,-133.5</points>
<intersection>29 1</intersection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-133.5,28.5,-133</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-133.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32,-134,32,-133.5</points>
<connection>
<GID>135</GID>
<name>IN_3</name></connection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-133.5,32,-133.5</points>
<intersection>28.5 0</intersection>
<intersection>32 1</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-43.5,-19.5,-35.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-93,-35.5,-93,-27.5</points>
<connection>
<GID>174</GID>
<name>OUT_3</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-93,-35.5,-19.5,-35.5</points>
<intersection>-93 1</intersection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-93,-27.5,-91.5,-27.5</points>
<intersection>-93 1</intersection>
<intersection>-91.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-91.5,-27.5,-91.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_4</name></connection>
<intersection>-27.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-43.5,-29.5,-35.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-95,-35.5,-95,-18.5</points>
<connection>
<GID>174</GID>
<name>OUT_1</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-18.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-95,-35.5,-29.5,-35.5</points>
<intersection>-95 1</intersection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-95,-18.5,-93.5,-18.5</points>
<intersection>-95 1</intersection>
<intersection>-93.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-93.5,-18.5,-93.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_6</name></connection>
<intersection>-18.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-43.5,-24.5,-35.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-94,-35.5,-94,-21.5</points>
<connection>
<GID>174</GID>
<name>OUT_2</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-21.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-94,-35.5,-24.5,-35.5</points>
<intersection>-94 1</intersection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-94,-21.5,-92.5,-21.5</points>
<intersection>-94 1</intersection>
<intersection>-92.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-92.5,-21.5,-92.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_5</name></connection>
<intersection>-21.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-43.5,-14.5,-35.5</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-77.5,-35.5,-77.5,-17</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-17 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-35.5,-14.5,-35.5</points>
<intersection>-77.5 1</intersection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-90.5,-17,-77.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_3</name></connection>
<intersection>-77.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-43.5,-9.5,-35.5</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-76.5,-35.5,-76.5,-17</points>
<connection>
<GID>175</GID>
<name>OUT_1</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-17 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-76.5,-35.5,-9.5,-35.5</points>
<intersection>-76.5 1</intersection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-89.5,-17,-76.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_2</name></connection>
<intersection>-76.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-43.5,-4.5,-35.5</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-75.5,-35.5,-75.5,-17</points>
<connection>
<GID>175</GID>
<name>OUT_2</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-17 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-75.5,-35.5,-4.5,-35.5</points>
<intersection>-75.5 1</intersection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-88.5,-17,-75.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>-75.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-43.5,0.5,-35.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-74.5,-35.5,-74.5,-17</points>
<connection>
<GID>175</GID>
<name>OUT_3</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-17 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-74.5,-35.5,0.5,-35.5</points>
<intersection>-74.5 1</intersection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-87.5,-17,-74.5,-17</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-74.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-134,30.5,-133</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-134 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30,-134,30.5,-134</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-21,18.5,-21</points>
<connection>
<GID>198</GID>
<name>carry_in</name></connection>
<connection>
<GID>199</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-133.5,29.5,-133</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-133.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,-134,31,-133.5</points>
<connection>
<GID>135</GID>
<name>IN_2</name></connection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-133.5,31,-133.5</points>
<intersection>29.5 0</intersection>
<intersection>31 1</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-43.5,-32.5,-34.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>28,-34.5,28,-26</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-32.5,-34.5,28,-34.5</points>
<intersection>-32.5 0</intersection>
<intersection>28 1</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-34.5,27,-26</points>
<connection>
<GID>199</GID>
<name>OUT_1</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-27.5,-43.5,-27.5,-34.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-34.5,27,-34.5</points>
<intersection>-27.5 1</intersection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-43.5,-22.5,-34.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26,-34.5,26,-26</points>
<connection>
<GID>199</GID>
<name>OUT_2</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-22.5,-34.5,26,-34.5</points>
<intersection>-22.5 0</intersection>
<intersection>26 1</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,-43.5,-17.5,-34.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25,-34.5,25,-26</points>
<connection>
<GID>199</GID>
<name>OUT_3</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-17.5,-34.5,25,-34.5</points>
<intersection>-17.5 0</intersection>
<intersection>25 1</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-43.5,-12.5,-34.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>9.5,-34.5,9.5,-26</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-34.5,9.5,-34.5</points>
<intersection>-12.5 0</intersection>
<intersection>9.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-43.5,-7.5,-34.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8.5,-34.5,8.5,-26</points>
<connection>
<GID>198</GID>
<name>OUT_1</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-34.5,8.5,-34.5</points>
<intersection>-7.5 0</intersection>
<intersection>8.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-43.5,-2.5,-34.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>7.5,-34.5,7.5,-26</points>
<connection>
<GID>198</GID>
<name>OUT_2</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2.5,-34.5,7.5,-34.5</points>
<intersection>-2.5 0</intersection>
<intersection>7.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-43.5,2.5,-34.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6.5,-34.5,6.5,-26</points>
<connection>
<GID>198</GID>
<name>OUT_3</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-34.5,6.5,-34.5</points>
<intersection>2.5 0</intersection>
<intersection>6.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-32,-15,-25</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-33.5,-39.5,-33.5,-32</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-32,-15,-32</points>
<intersection>-33.5 1</intersection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-32,-16,-25</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-28.5,-39.5,-28.5,-32</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-32,-16,-32</points>
<intersection>-28.5 1</intersection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-32,-17,-25</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-23.5,-39.5,-23.5,-32</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-32,-17,-32</points>
<intersection>-23.5 1</intersection>
<intersection>-17 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,-32,-18,-25</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-18.5,-39.5,-18.5,-32</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-18.5,-32,-18,-32</points>
<intersection>-18.5 1</intersection>
<intersection>-18 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,-32,-19,-25</points>
<connection>
<GID>60</GID>
<name>IN_4</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-13.5,-39.5,-13.5,-32</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-19,-32,-13.5,-32</points>
<intersection>-19 0</intersection>
<intersection>-13.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-32,-20,-25</points>
<connection>
<GID>60</GID>
<name>IN_5</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-8.5,-39.5,-8.5,-32</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-20,-32,-8.5,-32</points>
<intersection>-20 0</intersection>
<intersection>-8.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-32,-21,-25</points>
<connection>
<GID>60</GID>
<name>IN_6</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-3.5,-39.5,-3.5,-32</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-21,-32,-3.5,-32</points>
<intersection>-21 0</intersection>
<intersection>-3.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-32,-22,-25</points>
<connection>
<GID>60</GID>
<name>IN_7</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>1.5,-39.5,1.5,-32</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-22,-32,1.5,-32</points>
<intersection>-22 0</intersection>
<intersection>1.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-137,35,-137</points>
<connection>
<GID>135</GID>
<name>load</name></connection>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-93.5,56,-93</points>
<connection>
<GID>295</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,-94,53,-93.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53,-93.5,56,-93.5</points>
<intersection>53 1</intersection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-132,-15,-96,-15</points>
<connection>
<GID>209</GID>
<name>ENABLE_0</name></connection>
<intersection>-132 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>-132,-123.5,-132,-15</points>
<intersection>-123.5 2</intersection>
<intersection>-15 0</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-132,-123.5,31.5,-123.5</points>
<intersection>-132 1</intersection>
<intersection>31.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>31.5,-123.5,31.5,-122</points>
<connection>
<GID>132</GID>
<name>OUT_3</name></connection>
<intersection>-123.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-93.5,53,-93</points>
<connection>
<GID>295</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56,-94,56,-93.5</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53,-93.5,56,-93.5</points>
<intersection>53 0</intersection>
<intersection>56 1</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-93.5,55,-93</points>
<connection>
<GID>295</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>54,-94,54,-93.5</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-93.5,55,-93.5</points>
<intersection>54 1</intersection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-93.5,54,-93</points>
<connection>
<GID>295</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>55,-94,55,-93.5</points>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-93.5,55,-93.5</points>
<intersection>54 0</intersection>
<intersection>55 1</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-97,59,-97</points>
<connection>
<GID>138</GID>
<name>load</name></connection>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-113.5,56,-113</points>
<connection>
<GID>296</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-113 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52,-116,52,-113</points>
<intersection>-116 3</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52,-113,56,-113</points>
<intersection>52 1</intersection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,-116,53,-116</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>52 1</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-24,91.5,29.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>-24 5</intersection>
<intersection>29.5 9</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>91.5,-24,93.5,-24</points>
<connection>
<GID>231</GID>
<name>ENABLE_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>90.5,29.5,91.5,29.5</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-9,91.5,30.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>-9 5</intersection>
<intersection>30.5 9</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>91.5,-9,93.5,-9</points>
<connection>
<GID>230</GID>
<name>ENABLE_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>90.5,30.5,91.5,30.5</points>
<connection>
<GID>238</GID>
<name>OUT_1</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,6,91.5,31.5</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>6 5</intersection>
<intersection>31.5 9</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>91.5,6,93.5,6</points>
<connection>
<GID>229</GID>
<name>ENABLE_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>90.5,31.5,91.5,31.5</points>
<connection>
<GID>238</GID>
<name>OUT_2</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,21,91.5,32.5</points>
<connection>
<GID>243</GID>
<name>IN_3</name></connection>
<intersection>21 5</intersection>
<intersection>32.5 9</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>91.5,21,93.5,21</points>
<connection>
<GID>232</GID>
<name>ENABLE_0</name></connection>
<intersection>91.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>90.5,32.5,91.5,32.5</points>
<connection>
<GID>238</GID>
<name>OUT_3</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,7,117.5,7</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<connection>
<GID>246</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-8,117.5,-8</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<connection>
<GID>247</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,4.5,95.5,4.5</points>
<connection>
<GID>229</GID>
<name>OUT_7</name></connection>
<connection>
<GID>240</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-1.5,95.5,-1.5</points>
<connection>
<GID>229</GID>
<name>OUT_1</name></connection>
<connection>
<GID>240</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,0.5,95.5,0.5</points>
<connection>
<GID>229</GID>
<name>OUT_3</name></connection>
<connection>
<GID>240</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-0.5,95.5,-0.5</points>
<connection>
<GID>229</GID>
<name>OUT_2</name></connection>
<connection>
<GID>240</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-2.5,95.5,-2.5</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,3.5,95.5,3.5</points>
<connection>
<GID>229</GID>
<name>OUT_6</name></connection>
<connection>
<GID>240</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,1.5,95.5,1.5</points>
<connection>
<GID>229</GID>
<name>OUT_4</name></connection>
<connection>
<GID>240</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,2.5,95.5,2.5</points>
<connection>
<GID>229</GID>
<name>OUT_5</name></connection>
<connection>
<GID>240</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-17.5,95.5,-17.5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<connection>
<GID>241</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-15.5,95.5,-15.5</points>
<connection>
<GID>230</GID>
<name>OUT_2</name></connection>
<connection>
<GID>241</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-16.5,95.5,-16.5</points>
<connection>
<GID>230</GID>
<name>OUT_1</name></connection>
<connection>
<GID>241</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-14.5,95.5,-14.5</points>
<connection>
<GID>230</GID>
<name>OUT_3</name></connection>
<connection>
<GID>241</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-13.5,95.5,-13.5</points>
<connection>
<GID>230</GID>
<name>OUT_4</name></connection>
<connection>
<GID>241</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-12.5,95.5,-12.5</points>
<connection>
<GID>230</GID>
<name>OUT_5</name></connection>
<connection>
<GID>241</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-10.5,95.5,-10.5</points>
<connection>
<GID>230</GID>
<name>OUT_7</name></connection>
<connection>
<GID>241</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-11.5,95.5,-11.5</points>
<connection>
<GID>230</GID>
<name>OUT_6</name></connection>
<connection>
<GID>241</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,13.5,95.5,13.5</points>
<connection>
<GID>232</GID>
<name>OUT_1</name></connection>
<connection>
<GID>239</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,15.5,95.5,15.5</points>
<connection>
<GID>232</GID>
<name>OUT_3</name></connection>
<connection>
<GID>239</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,16.5,95.5,16.5</points>
<connection>
<GID>232</GID>
<name>OUT_4</name></connection>
<connection>
<GID>239</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,12.5,95.5,12.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<connection>
<GID>239</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,14.5,95.5,14.5</points>
<connection>
<GID>232</GID>
<name>OUT_2</name></connection>
<connection>
<GID>239</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,17.5,95.5,17.5</points>
<connection>
<GID>232</GID>
<name>OUT_5</name></connection>
<connection>
<GID>239</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,18.5,95.5,18.5</points>
<connection>
<GID>232</GID>
<name>OUT_6</name></connection>
<connection>
<GID>239</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,19.5,95.5,19.5</points>
<connection>
<GID>232</GID>
<name>OUT_7</name></connection>
<connection>
<GID>239</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-26.5,95.5,-26.5</points>
<connection>
<GID>231</GID>
<name>OUT_6</name></connection>
<connection>
<GID>242</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-31.5,95.5,-31.5</points>
<connection>
<GID>231</GID>
<name>OUT_1</name></connection>
<connection>
<GID>242</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-28.5,95.5,-28.5</points>
<connection>
<GID>231</GID>
<name>OUT_4</name></connection>
<connection>
<GID>242</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-25.5,95.5,-25.5</points>
<connection>
<GID>231</GID>
<name>OUT_7</name></connection>
<connection>
<GID>242</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-29.5,95.5,-29.5</points>
<connection>
<GID>231</GID>
<name>OUT_3</name></connection>
<connection>
<GID>242</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-32.5,95.5,-32.5</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<connection>
<GID>242</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-30.5,95.5,-30.5</points>
<connection>
<GID>231</GID>
<name>OUT_2</name></connection>
<connection>
<GID>242</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-27.5,95.5,-27.5</points>
<connection>
<GID>231</GID>
<name>OUT_5</name></connection>
<connection>
<GID>242</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-144,93.5,34</points>
<connection>
<GID>243</GID>
<name>ENABLE_0</name></connection>
<intersection>-144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-144,93.5,-144</points>
<intersection>29.5 2</intersection>
<intersection>93.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>29.5,-144,29.5,-142</points>
<intersection>-144 1</intersection>
<intersection>-142 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29.5,-142,31,-142</points>
<connection>
<GID>135</GID>
<name>OUT_2</name></connection>
<intersection>29.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-23.5,95.5,29.5</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-23.5,98.5,-23.5</points>
<connection>
<GID>242</GID>
<name>load</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-8.5,95.5,30.5</points>
<connection>
<GID>243</GID>
<name>OUT_1</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-8.5,98.5,-8.5</points>
<connection>
<GID>241</GID>
<name>load</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,6.5,95.5,31.5</points>
<connection>
<GID>243</GID>
<name>OUT_2</name></connection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95.5,6.5,98.5,6.5</points>
<connection>
<GID>240</GID>
<name>load</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,21.5,95.5,32.5</points>
<connection>
<GID>243</GID>
<name>OUT_3</name></connection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95.5,21.5,98.5,21.5</points>
<connection>
<GID>239</GID>
<name>load</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-115,53,-113.5</points>
<connection>
<GID>296</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-115 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56,-116,56,-115</points>
<connection>
<GID>140</GID>
<name>IN_3</name></connection>
<intersection>-115 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53,-115,56,-115</points>
<intersection>53 0</intersection>
<intersection>56 1</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,19.5</points>
<intersection>-11 4</intersection>
<intersection>4 1</intersection>
<intersection>19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>248</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,19.5,104.5,19.5</points>
<connection>
<GID>239</GID>
<name>OUT_7</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>259</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,4.5</points>
<intersection>-13 4</intersection>
<intersection>2 1</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>248</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,4.5,104.5,4.5</points>
<connection>
<GID>240</GID>
<name>OUT_7</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>259</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-15,104.5,0</points>
<intersection>-15 3</intersection>
<intersection>-10.5 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-10.5,104.5,-10.5</points>
<connection>
<GID>241</GID>
<name>OUT_7</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-25.5,104.5,-2</points>
<intersection>-25.5 2</intersection>
<intersection>-17 3</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-25.5,104.5,-25.5</points>
<connection>
<GID>242</GID>
<name>OUT_7</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,18.5</points>
<intersection>-11 4</intersection>
<intersection>4 1</intersection>
<intersection>18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>249</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,18.5,104.5,18.5</points>
<connection>
<GID>239</GID>
<name>OUT_6</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>263</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,3.5</points>
<intersection>-13 4</intersection>
<intersection>2 1</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>249</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,3.5,104.5,3.5</points>
<connection>
<GID>240</GID>
<name>OUT_6</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>263</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<intersection>104.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>104.5,-15,104.5,0</points>
<intersection>-15 5</intersection>
<intersection>-11.5 4</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>103.5,-11.5,104.5,-11.5</points>
<connection>
<GID>241</GID>
<name>OUT_6</name></connection>
<intersection>104.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>104.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-26.5,104.5,-2</points>
<intersection>-26.5 2</intersection>
<intersection>-17 3</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-26.5,104.5,-26.5</points>
<connection>
<GID>242</GID>
<name>OUT_6</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,1,113.5,5</points>
<intersection>1 3</intersection>
<intersection>5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>111.5,1,113.5,1</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>113.5,5,165.5,5</points>
<connection>
<GID>246</GID>
<name>IN_7</name></connection>
<connection>
<GID>225</GID>
<name>IN_7</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,1,113.5,4</points>
<intersection>1 2</intersection>
<intersection>4 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,1,113.5,1</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>113.5,4,165.5,4</points>
<connection>
<GID>246</GID>
<name>IN_6</name></connection>
<connection>
<GID>225</GID>
<name>IN_6</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,6,109.5,28.5</points>
<connection>
<GID>258</GID>
<name>SEL_0</name></connection>
<connection>
<GID>257</GID>
<name>SEL_0</name></connection>
<connection>
<GID>256</GID>
<name>SEL_0</name></connection>
<connection>
<GID>255</GID>
<name>SEL_0</name></connection>
<connection>
<GID>254</GID>
<name>SEL_0</name></connection>
<connection>
<GID>253</GID>
<name>SEL_0</name></connection>
<connection>
<GID>249</GID>
<name>SEL_0</name></connection>
<connection>
<GID>248</GID>
<name>SEL_0</name></connection>
<intersection>28.5 145</intersection></vsegment>
<hsegment>
<ID>145</ID>
<points>106,28.5,109.5,28.5</points>
<connection>
<GID>244</GID>
<name>N_in1</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,6,108.5,31.5</points>
<connection>
<GID>258</GID>
<name>SEL_1</name></connection>
<connection>
<GID>257</GID>
<name>SEL_1</name></connection>
<connection>
<GID>256</GID>
<name>SEL_1</name></connection>
<connection>
<GID>255</GID>
<name>SEL_1</name></connection>
<connection>
<GID>254</GID>
<name>SEL_1</name></connection>
<connection>
<GID>253</GID>
<name>SEL_1</name></connection>
<connection>
<GID>249</GID>
<name>SEL_1</name></connection>
<connection>
<GID>248</GID>
<name>SEL_1</name></connection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,31.5,108.5,31.5</points>
<connection>
<GID>235</GID>
<name>N_in1</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,17.5</points>
<intersection>-11 7</intersection>
<intersection>4 1</intersection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>253</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,17.5,104.5,17.5</points>
<connection>
<GID>239</GID>
<name>OUT_5</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>264</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,2.5</points>
<intersection>-13 7</intersection>
<intersection>2 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>253</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,2.5,104.5,2.5</points>
<connection>
<GID>240</GID>
<name>OUT_5</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>264</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-15,104.5,0</points>
<intersection>-15 3</intersection>
<intersection>-12.5 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-12.5,104.5,-12.5</points>
<connection>
<GID>241</GID>
<name>OUT_5</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-27.5,104.5,-2</points>
<intersection>-27.5 2</intersection>
<intersection>-17 3</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-27.5,104.5,-27.5</points>
<connection>
<GID>242</GID>
<name>OUT_5</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,1,113.5,3</points>
<intersection>1 2</intersection>
<intersection>3 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,1,113.5,1</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>113.5,3,165.5,3</points>
<connection>
<GID>246</GID>
<name>IN_5</name></connection>
<connection>
<GID>225</GID>
<name>IN_5</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,16.5</points>
<intersection>-11 4</intersection>
<intersection>4 1</intersection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>254</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,16.5,104.5,16.5</points>
<connection>
<GID>239</GID>
<name>OUT_4</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>265</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,2</points>
<intersection>-13 3</intersection>
<intersection>1.5 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>254</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,1.5,104.5,1.5</points>
<connection>
<GID>240</GID>
<name>OUT_4</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>265</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-15,104.5,0</points>
<intersection>-15 3</intersection>
<intersection>-13.5 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-13.5,104.5,-13.5</points>
<connection>
<GID>241</GID>
<name>OUT_4</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-28.5,104.5,-2</points>
<intersection>-28.5 2</intersection>
<intersection>-17 3</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-28.5,104.5,-28.5</points>
<connection>
<GID>242</GID>
<name>OUT_4</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>111.5,5.5,113.5,5.5</points>
<intersection>111.5 4</intersection>
<intersection>113.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>111.5,1,111.5,5.5</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<intersection>5.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>113.5,2,113.5,5.5</points>
<intersection>2 6</intersection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>113.5,2,165.5,2</points>
<connection>
<GID>246</GID>
<name>IN_4</name></connection>
<connection>
<GID>225</GID>
<name>IN_4</name></connection>
<intersection>113.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,15.5</points>
<intersection>-11 4</intersection>
<intersection>4 1</intersection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>255</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,15.5,104.5,15.5</points>
<connection>
<GID>239</GID>
<name>OUT_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>266</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,2</points>
<intersection>-13 3</intersection>
<intersection>0.5 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>255</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,0.5,104.5,0.5</points>
<connection>
<GID>240</GID>
<name>OUT_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>266</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-15,104.5,0</points>
<intersection>-15 3</intersection>
<intersection>-14.5 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-14.5,104.5,-14.5</points>
<connection>
<GID>241</GID>
<name>OUT_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-29.5,104.5,-2</points>
<intersection>-29.5 2</intersection>
<intersection>-17 3</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-29.5,104.5,-29.5</points>
<connection>
<GID>242</GID>
<name>OUT_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111.5,5.5,113.5,5.5</points>
<intersection>111.5 4</intersection>
<intersection>113.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>111.5,1,111.5,5.5</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<intersection>5.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>113.5,1.5,113.5,5.5</points>
<intersection>1.5 6</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>113.5,1.5,114.5,1.5</points>
<intersection>113.5 5</intersection>
<intersection>114.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>114.5,1,114.5,1.5</points>
<connection>
<GID>246</GID>
<name>IN_3</name></connection>
<intersection>1 10</intersection>
<intersection>1.5 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>114.5,1,165.5,1</points>
<connection>
<GID>225</GID>
<name>IN_3</name></connection>
<intersection>114.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,14.5</points>
<intersection>-11 4</intersection>
<intersection>4 2</intersection>
<intersection>14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,14.5,104.5,14.5</points>
<connection>
<GID>239</GID>
<name>OUT_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>256</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>267</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,2</points>
<intersection>-13 3</intersection>
<intersection>-0.5 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-0.5,104.5,-0.5</points>
<connection>
<GID>240</GID>
<name>OUT_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>256</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>267</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-15.5,104.5,0</points>
<intersection>-15.5 1</intersection>
<intersection>-15 3</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-15.5,104.5,-15.5</points>
<connection>
<GID>241</GID>
<name>OUT_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-30.5,104.5,-2</points>
<intersection>-30.5 1</intersection>
<intersection>-17 3</intersection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-30.5,104.5,-30.5</points>
<connection>
<GID>242</GID>
<name>OUT_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,0,113.5,1</points>
<intersection>0 5</intersection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,1,113.5,1</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>113.5,0,165.5,0</points>
<connection>
<GID>246</GID>
<name>IN_2</name></connection>
<connection>
<GID>225</GID>
<name>IN_2</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,13.5</points>
<intersection>-11 7</intersection>
<intersection>4 2</intersection>
<intersection>13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,13.5,104.5,13.5</points>
<connection>
<GID>239</GID>
<name>OUT_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>257</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>268</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,2</points>
<intersection>-13 1</intersection>
<intersection>-1.5 5</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>268</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>257</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103.5,-1.5,104.5,-1.5</points>
<connection>
<GID>240</GID>
<name>OUT_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-16.5,104.5,0</points>
<intersection>-16.5 1</intersection>
<intersection>-15 3</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-16.5,104.5,-16.5</points>
<connection>
<GID>241</GID>
<name>OUT_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-31.5,104.5,-2</points>
<intersection>-31.5 1</intersection>
<intersection>-17 3</intersection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-31.5,104.5,-31.5</points>
<connection>
<GID>242</GID>
<name>OUT_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-1,113,1</points>
<intersection>-1 5</intersection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,1,113,1</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>113,-1,165.5,-1</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-2,113.5,1</points>
<intersection>-2 5</intersection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,1,113.5,1</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>113.5,-2,165.5,-2</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-11,104.5,12.5</points>
<intersection>-11 8</intersection>
<intersection>4 2</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,12.5,104.5,12.5</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,4,105.5,4</points>
<connection>
<GID>258</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>104.5,-11,105.5,-11</points>
<connection>
<GID>269</GID>
<name>IN_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-13,104.5,2</points>
<intersection>-13 3</intersection>
<intersection>-2.5 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-2.5,104.5,-2.5</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,2,105.5,2</points>
<connection>
<GID>258</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-13,105.5,-13</points>
<connection>
<GID>269</GID>
<name>IN_2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-17.5,104.5,0</points>
<intersection>-17.5 1</intersection>
<intersection>-15 3</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-17.5,104.5,-17.5</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,0,105.5,0</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-15,105.5,-15</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-32.5,104.5,-2</points>
<intersection>-32.5 1</intersection>
<intersection>-17 3</intersection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-32.5,104.5,-32.5</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-2,105.5,-2</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-17,105.5,-17</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-9,108.5,31.5</points>
<connection>
<GID>269</GID>
<name>SEL_1</name></connection>
<connection>
<GID>268</GID>
<name>SEL_1</name></connection>
<connection>
<GID>267</GID>
<name>SEL_1</name></connection>
<connection>
<GID>266</GID>
<name>SEL_1</name></connection>
<connection>
<GID>265</GID>
<name>SEL_1</name></connection>
<connection>
<GID>264</GID>
<name>SEL_1</name></connection>
<connection>
<GID>263</GID>
<name>SEL_1</name></connection>
<connection>
<GID>259</GID>
<name>SEL_1</name></connection>
<intersection>31.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>108.5,31.5,111,31.5</points>
<connection>
<GID>279</GID>
<name>N_in0</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-9,109.5,28.5</points>
<connection>
<GID>269</GID>
<name>SEL_0</name></connection>
<connection>
<GID>268</GID>
<name>SEL_0</name></connection>
<connection>
<GID>267</GID>
<name>SEL_0</name></connection>
<connection>
<GID>266</GID>
<name>SEL_0</name></connection>
<connection>
<GID>265</GID>
<name>SEL_0</name></connection>
<connection>
<GID>264</GID>
<name>SEL_0</name></connection>
<connection>
<GID>263</GID>
<name>SEL_0</name></connection>
<connection>
<GID>259</GID>
<name>SEL_0</name></connection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,28.5,111,28.5</points>
<connection>
<GID>281</GID>
<name>N_in0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-14,113.5,-10</points>
<intersection>-14 2</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-10,114.5,-10</points>
<connection>
<GID>247</GID>
<name>IN_7</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-14,113.5,-14</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-14,113.5,-11</points>
<intersection>-14 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-11,114.5,-11</points>
<connection>
<GID>247</GID>
<name>IN_6</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-14,113.5,-14</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-14,113.5,-12</points>
<intersection>-14 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-12,114.5,-12</points>
<connection>
<GID>247</GID>
<name>IN_5</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-14,113.5,-14</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-14,113.5,-13</points>
<intersection>-14 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-13,114.5,-13</points>
<connection>
<GID>247</GID>
<name>IN_4</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-14,113.5,-14</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111.5,-14,114.5,-14</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<connection>
<GID>247</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-15,113.5,-14</points>
<intersection>-15 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-15,114.5,-15</points>
<connection>
<GID>247</GID>
<name>IN_2</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-14,113.5,-14</points>
<connection>
<GID>267</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-16,113.5,-14</points>
<intersection>-16 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-16,114.5,-16</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-14,113.5,-14</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-17,113.5,-14</points>
<intersection>-17 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-17,114.5,-17</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-14,113.5,-14</points>
<connection>
<GID>269</GID>
<name>OUT</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-114.5,54.5,-113.5</points>
<intersection>-114.5 2</intersection>
<intersection>-113.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>54,-116,54,-114.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>-114.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-114.5,54.5,-114.5</points>
<intersection>54 1</intersection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54.5,-113.5,55,-113.5</points>
<connection>
<GID>296</GID>
<name>DATA_OUT_1</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-97,143,-97</points>
<connection>
<GID>319</GID>
<name>carry_out</name></connection>
<connection>
<GID>320</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-94,156,-91.5</points>
<connection>
<GID>319</GID>
<name>IN_B_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>158,-91.5,158,-17</points>
<intersection>-91.5 2</intersection>
<intersection>-17 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117,-91.5,158,-91.5</points>
<intersection>117 4</intersection>
<intersection>156 0</intersection>
<intersection>158 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>117,-95,117,-91.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>122.5,-17,158,-17</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>158 1</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-94,155,-16</points>
<connection>
<GID>319</GID>
<name>IN_B_1</name></connection>
<intersection>-90.5 2</intersection>
<intersection>-16 18</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117,-90.5,155,-90.5</points>
<intersection>117 3</intersection>
<intersection>155 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-95,117,-90.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>122.5,-16,155,-16</points>
<connection>
<GID>247</GID>
<name>OUT_1</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-94,154,-91.5</points>
<connection>
<GID>319</GID>
<name>IN_B_2</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>152,-91.5,152,-15</points>
<intersection>-91.5 2</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117,-91.5,154,-91.5</points>
<intersection>117 5</intersection>
<intersection>152 1</intersection>
<intersection>154 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>117,-95,117,-91.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>122.5,-15,152,-15</points>
<connection>
<GID>247</GID>
<name>OUT_2</name></connection>
<intersection>152 1</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-94,153,-91.5</points>
<connection>
<GID>319</GID>
<name>IN_B_3</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>149,-91.5,149,-14</points>
<intersection>-91.5 2</intersection>
<intersection>-14 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117,-91.5,153,-91.5</points>
<intersection>117 4</intersection>
<intersection>149 1</intersection>
<intersection>153 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>117,-95,117,-91.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>122.5,-14,149,-14</points>
<connection>
<GID>247</GID>
<name>OUT_3</name></connection>
<intersection>149 1</intersection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-94,149,-93</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,149,-93</points>
<intersection>115 4</intersection>
<intersection>122.5 15</intersection>
<intersection>149 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>330</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>122.5,-93,122.5,-2</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-94,148,-93</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,148,-93</points>
<intersection>115 4</intersection>
<intersection>122.5 15</intersection>
<intersection>148 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>122.5,-93,122.5,-1</points>
<connection>
<GID>246</GID>
<name>OUT_1</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-94,147,-93</points>
<connection>
<GID>319</GID>
<name>IN_2</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,147,-93</points>
<intersection>115 5</intersection>
<intersection>122.5 16</intersection>
<intersection>147 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>122.5,-93,122.5,0</points>
<connection>
<GID>246</GID>
<name>OUT_2</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-94,146,-93</points>
<connection>
<GID>319</GID>
<name>IN_3</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,146,-93</points>
<intersection>115 4</intersection>
<intersection>122.5 15</intersection>
<intersection>146 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>122.5,-93,122.5,1</points>
<connection>
<GID>246</GID>
<name>OUT_3</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-94,133,-93</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,133,-93</points>
<intersection>115 4</intersection>
<intersection>122.5 15</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>122.5,-93,122.5,2</points>
<connection>
<GID>246</GID>
<name>OUT_4</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-94,132,-93</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,132,-93</points>
<intersection>115 10</intersection>
<intersection>122.5 21</intersection>
<intersection>132 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>122.5,-93,122.5,3</points>
<connection>
<GID>246</GID>
<name>OUT_5</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-94,131,-93</points>
<connection>
<GID>320</GID>
<name>IN_2</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,131,-93</points>
<intersection>115 8</intersection>
<intersection>122.5 11</intersection>
<intersection>131 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>122.5,-93,122.5,4</points>
<connection>
<GID>246</GID>
<name>OUT_6</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-94,130,-93</points>
<connection>
<GID>320</GID>
<name>IN_3</name></connection>
<intersection>-93 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>115,-95,115,-93</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-93,130,-93</points>
<intersection>115 1</intersection>
<intersection>122.5 21</intersection>
<intersection>130 0</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>122.5,-93,122.5,5</points>
<connection>
<GID>246</GID>
<name>OUT_7</name></connection>
<intersection>-93 2</intersection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-94,137,-10</points>
<connection>
<GID>320</GID>
<name>IN_B_3</name></connection>
<intersection>-90.5 3</intersection>
<intersection>-10 19</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>117,-90.5,137,-90.5</points>
<intersection>117 4</intersection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>117,-95,117,-90.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>-90.5 3</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>122.5,-10,137,-10</points>
<connection>
<GID>247</GID>
<name>OUT_7</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-95,117,-91.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>-94 10</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117,-91.5,140,-91.5</points>
<intersection>117 0</intersection>
<intersection>140 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>140,-91.5,140,-11</points>
<intersection>-91.5 2</intersection>
<intersection>-11 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>122.5,-11,140,-11</points>
<connection>
<GID>247</GID>
<name>OUT_6</name></connection>
<intersection>140 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>117,-94,138,-94</points>
<connection>
<GID>320</GID>
<name>IN_B_2</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-94,139,-91.5</points>
<connection>
<GID>320</GID>
<name>IN_B_1</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>143,-91.5,143,-12</points>
<intersection>-91.5 2</intersection>
<intersection>-12 13</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117,-91.5,143,-91.5</points>
<intersection>117 12</intersection>
<intersection>139 0</intersection>
<intersection>143 1</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>117,-95,117,-91.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>122.5,-12,143,-12</points>
<connection>
<GID>247</GID>
<name>OUT_5</name></connection>
<intersection>143 1</intersection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-95,117,-91.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>146,-91.5,146,-13</points>
<intersection>-91.5 2</intersection>
<intersection>-13 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117,-91.5,146,-91.5</points>
<intersection>117 0</intersection>
<intersection>140 7</intersection>
<intersection>146 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>140,-94,140,-91.5</points>
<connection>
<GID>320</GID>
<name>IN_B_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>122.5,-13,146,-13</points>
<connection>
<GID>247</GID>
<name>OUT_4</name></connection>
<intersection>146 1</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-104,146.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_7</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>152.5,-103,152.5,-102</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>146.5,-103,152.5,-103</points>
<intersection>146.5 0</intersection>
<intersection>152.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-104,145.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_6</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>151.5,-103,151.5,-102</points>
<connection>
<GID>319</GID>
<name>OUT_1</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>145.5,-103,151.5,-103</points>
<intersection>145.5 0</intersection>
<intersection>151.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-104,144.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_5</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>150.5,-103,150.5,-102</points>
<connection>
<GID>319</GID>
<name>OUT_2</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>144.5,-103,150.5,-103</points>
<intersection>144.5 0</intersection>
<intersection>150.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,-104,143.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_4</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>149.5,-103,149.5,-102</points>
<connection>
<GID>319</GID>
<name>OUT_3</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-103,149.5,-103</points>
<intersection>143.5 0</intersection>
<intersection>149.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-104,142.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_3</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>136.5,-103,136.5,-102</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>136.5,-103,142.5,-103</points>
<intersection>136.5 1</intersection>
<intersection>142.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-104,141.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_2</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>135.5,-103,135.5,-102</points>
<connection>
<GID>320</GID>
<name>OUT_1</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>135.5,-103,141.5,-103</points>
<intersection>135.5 1</intersection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-104,140.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>134.5,-103,134.5,-102</points>
<connection>
<GID>320</GID>
<name>OUT_2</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134.5,-103,140.5,-103</points>
<intersection>134.5 1</intersection>
<intersection>140.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-104,139.5,-103</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>133.5,-103,133.5,-102</points>
<connection>
<GID>320</GID>
<name>OUT_3</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>133.5,-103,139.5,-103</points>
<intersection>133.5 1</intersection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-104,112.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-103,116,-103</points>
<intersection>112.5 0</intersection>
<intersection>116 1</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<intersection>-103 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>113.5,-103,116,-103</points>
<intersection>113.5 10</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>113.5,-104,113.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_1</name></connection>
<intersection>-103 9</intersection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-104,114.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_2</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-103,116,-103</points>
<intersection>114.5 0</intersection>
<intersection>116 1</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-104,115.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_3</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-103,116,-103</points>
<intersection>115.5 0</intersection>
<intersection>116 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>-103 2</intersection></vsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-104,116.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_4</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>116,-103,116.5,-103</points>
<intersection>116 3</intersection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>-103 2</intersection></vsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-104,117.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_5</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>116,-103,117.5,-103</points>
<intersection>116 1</intersection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-104,118.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_6</name></connection>
<intersection>-103 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>116,-103,118.5,-103</points>
<intersection>116 1</intersection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-104,119.5,-103</points>
<connection>
<GID>324</GID>
<name>IN_7</name></connection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>116,-103,119.5,-103</points>
<intersection>116 3</intersection>
<intersection>119.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116,-103,116,-101</points>
<connection>
<GID>330</GID>
<name>OUT</name></connection>
<intersection>-103 2</intersection></vsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>112.5,-108,139.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>113.5,-108,140.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<connection>
<GID>324</GID>
<name>OUT_1</name></connection>
<connection>
<GID>321</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>114.5,-108,141.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_2</name></connection>
<connection>
<GID>324</GID>
<name>OUT_2</name></connection>
<connection>
<GID>321</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>115.5,-108,142.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_3</name></connection>
<connection>
<GID>324</GID>
<name>OUT_3</name></connection>
<connection>
<GID>321</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>116.5,-108,143.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_4</name></connection>
<connection>
<GID>324</GID>
<name>OUT_4</name></connection>
<connection>
<GID>321</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>117.5,-108,144.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_5</name></connection>
<connection>
<GID>324</GID>
<name>OUT_5</name></connection>
<connection>
<GID>321</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>118.5,-108,145.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_6</name></connection>
<connection>
<GID>324</GID>
<name>OUT_6</name></connection>
<connection>
<GID>321</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>119.5,-108,146.5,-108</points>
<connection>
<GID>332</GID>
<name>IN_7</name></connection>
<connection>
<GID>324</GID>
<name>OUT_7</name></connection>
<connection>
<GID>321</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-113,123.5,-112</points>
<connection>
<GID>333</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-112,130.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-113,126.5,-112</points>
<connection>
<GID>334</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>126.5,-112,131.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_1</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-113,129.5,-112</points>
<connection>
<GID>335</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-112,132.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-113,132.5,-112</points>
<connection>
<GID>336</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-112,133.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_3</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-113,135.5,-112</points>
<connection>
<GID>337</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134.5,-112,135.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_4</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-113,138.5,-112</points>
<connection>
<GID>338</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>135.5,-112,138.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_5</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-113,141.5,-112</points>
<connection>
<GID>339</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>136.5,-112,141.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_6</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-113,144.5,-112</points>
<connection>
<GID>340</GID>
<name>N_in3</name></connection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-112,144.5,-112</points>
<connection>
<GID>332</GID>
<name>OUT_7</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-106,148,-106</points>
<connection>
<GID>321</GID>
<name>ENABLE_0</name></connection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>125,-126,125,-106</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>-126 19</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>55,-126,125,-126</points>
<intersection>55 21</intersection>
<intersection>125 4</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>55,-126,55,-124</points>
<connection>
<GID>140</GID>
<name>OUT_2</name></connection>
<intersection>-126 19</intersection></vsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-125,139,-125</points>
<intersection>29.5 6</intersection>
<intersection>139 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>139,-125,139,-110</points>
<connection>
<GID>332</GID>
<name>ENABLE_0</name></connection>
<intersection>-125 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>29.5,-125,29.5,-122</points>
<connection>
<GID>132</GID>
<name>OUT_1</name></connection>
<intersection>-125 1</intersection></vsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-106,121,-106</points>
<connection>
<GID>324</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-109,-13.5,-102</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<connection>
<GID>344</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-109,-10,-84</points>
<intersection>-109 4</intersection>
<intersection>-84 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-10,-84,32,-84</points>
<intersection>-10 0</intersection>
<intersection>32 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-11.5,-109,-10,-109</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>32,-84,32,-83.5</points>
<connection>
<GID>121</GID>
<name>OUT_3</name></connection>
<intersection>-84 3</intersection></vsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-103.5,-12.5,-96</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>-103.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-103.5,32,-103.5</points>
<intersection>-12.5 0</intersection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-103.5,32,-102.5</points>
<connection>
<GID>124</GID>
<name>OUT_3</name></connection>
<intersection>-103.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-18,24.5,-14</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-107.5,-142,-107.5,-142</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<connection>
<GID>364</GID>
<name>CLK</name></connection></vsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-148.5,-108,-144</points>
<intersection>-148.5 5</intersection>
<intersection>-144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,-144,-107.5,-144</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-109,-148.5,-108,-148.5</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-118.5,-8,-84</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8,-84,31,-84</points>
<intersection>-8 0</intersection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-84,31,-83.5</points>
<connection>
<GID>121</GID>
<name>OUT_2</name></connection>
<intersection>-84 2</intersection></vsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-114,54,-113.5</points>
<connection>
<GID>296</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-114 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>55,-116,55,-114</points>
<connection>
<GID>140</GID>
<name>IN_2</name></connection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-114,55,-114</points>
<intersection>54 0</intersection>
<intersection>55 1</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-119,59,-117.5</points>
<connection>
<GID>140</GID>
<name>load</name></connection>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-164,6.5,-102</points>
<connection>
<GID>2</GID>
<name>load</name></connection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-102,56,-102</points>
<connection>
<GID>138</GID>
<name>OUT_3</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>1262.57,1845.1,3040.57,927.1</PageViewport>
<gate>
<ID>195</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>1284,709</position>
<output>
<ID>OUT_0</ID>224 </output>
<output>
<ID>OUT_1</ID>225 </output>
<output>
<ID>OUT_2</ID>386 </output>
<output>
<ID>OUT_3</ID>391 </output>
<output>
<ID>OUT_4</ID>392 </output>
<output>
<ID>OUT_5</ID>400 </output>
<output>
<ID>OUT_6</ID>403 </output>
<output>
<ID>OUT_7</ID>406 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_RAM_8x8</type>
<position>1323,682</position>
<input>
<ID>DATA_IN_0</ID>178 </input>
<input>
<ID>DATA_IN_1</ID>140 </input>
<input>
<ID>DATA_IN_2</ID>135 </input>
<input>
<ID>DATA_IN_3</ID>134 </input>
<input>
<ID>DATA_IN_4</ID>133 </input>
<input>
<ID>DATA_IN_5</ID>132 </input>
<input>
<ID>DATA_IN_6</ID>24 </input>
<input>
<ID>DATA_IN_7</ID>10 </input>
<output>
<ID>DATA_OUT_0</ID>178 </output>
<output>
<ID>DATA_OUT_1</ID>140 </output>
<output>
<ID>DATA_OUT_2</ID>135 </output>
<output>
<ID>DATA_OUT_3</ID>134 </output>
<output>
<ID>DATA_OUT_4</ID>133 </output>
<output>
<ID>DATA_OUT_5</ID>132 </output>
<output>
<ID>DATA_OUT_6</ID>24 </output>
<output>
<ID>DATA_OUT_7</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>8</ID>
<type>EE_VDD</type>
<position>666,-81.5</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>EE_VDD</type>
<position>673.5,-81.5</position>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>650,-92</position>
<gparam>LABEL_TEXT MSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>673,-91.5</position>
<gparam>LABEL_TEXT LSB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>673.5,-39</position>
<gparam>LABEL_TEXT BEN</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>695,-53.5</position>
<gparam>LABEL_TEXT COND + IRD</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_MUX_2x1</type>
<position>657,-84.5</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>34 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_OR2</type>
<position>666,-75.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_MUX_2x1</type>
<position>665,-84.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>35 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_MUX_2x1</type>
<position>672.5,-84.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>125 </input>
<output>
<ID>OUT</ID>56 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_MUX_2x1</type>
<position>650.5,-84.5</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>33 </output>
<input>
<ID>SEL_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_OR2</type>
<position>651.5,-76</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AE_OR3</type>
<position>666.5,-39.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<input>
<ID>IN_2</ID>129 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>49</ID>
<type>BA_ROM_4x4</type>
<position>695,-89.5</position>
<input>
<ID>ADDRESS_0</ID>56 </input>
<input>
<ID>ADDRESS_1</ID>35 </input>
<input>
<ID>ADDRESS_2</ID>34 </input>
<input>
<ID>ADDRESS_3</ID>33 </input>
<input>
<ID>ENABLE_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<gate>
<ID>50</ID>
<type>BA_ROM_4x4</type>
<position>694.5,-44</position>
<input>
<ID>ADDRESS_0</ID>56 </input>
<input>
<ID>ADDRESS_1</ID>35 </input>
<input>
<ID>ADDRESS_2</ID>34 </input>
<input>
<ID>ADDRESS_3</ID>33 </input>
<output>
<ID>DATA_OUT_0</ID>65 </output>
<output>
<ID>DATA_OUT_1</ID>55 </output>
<output>
<ID>DATA_OUT_2</ID>108 </output>
<output>
<ID>DATA_OUT_3</ID>82 </output>
<input>
<ID>ENABLE_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<gate>
<ID>51</ID>
<type>BA_ROM_4x4</type>
<position>694.5,-56.5</position>
<input>
<ID>ADDRESS_0</ID>56 </input>
<input>
<ID>ADDRESS_1</ID>35 </input>
<input>
<ID>ADDRESS_2</ID>34 </input>
<input>
<ID>ADDRESS_3</ID>33 </input>
<output>
<ID>DATA_OUT_0</ID>25 </output>
<output>
<ID>DATA_OUT_1</ID>67 </output>
<output>
<ID>DATA_OUT_3</ID>83 </output>
<input>
<ID>ENABLE_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>BA_ROM_4x4</type>
<position>694.5,-71.5</position>
<input>
<ID>ADDRESS_0</ID>56 </input>
<input>
<ID>ADDRESS_1</ID>35 </input>
<input>
<ID>ADDRESS_2</ID>34 </input>
<input>
<ID>ADDRESS_3</ID>33 </input>
<input>
<ID>ENABLE_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>693,-41</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>667,-69.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>EE_VDD</type>
<position>700.5,-44.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>EE_VDD</type>
<position>700.5,-57</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>59</ID>
<type>EE_VDD</type>
<position>700.5,-72</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>61</ID>
<type>EE_VDD</type>
<position>701,-90</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>63</ID>
<type>EE_VDD</type>
<position>724.5,-62.5</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>64</ID>
<type>EE_VDD</type>
<position>724.5,-80.5</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>65</ID>
<type>BA_ROM_4x4</type>
<position>718.5,-62</position>
<input>
<ID>ADDRESS_0</ID>56 </input>
<input>
<ID>ADDRESS_1</ID>35 </input>
<input>
<ID>ADDRESS_2</ID>34 </input>
<input>
<ID>ADDRESS_3</ID>33 </input>
<input>
<ID>ENABLE_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<gate>
<ID>66</ID>
<type>BA_ROM_4x4</type>
<position>718.5,-80</position>
<input>
<ID>ADDRESS_0</ID>56 </input>
<input>
<ID>ADDRESS_1</ID>35 </input>
<input>
<ID>ADDRESS_2</ID>34 </input>
<input>
<ID>ADDRESS_3</ID>33 </input>
<input>
<ID>ENABLE_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>650.5,-63</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>694.5,-82.5</position>
<gparam>LABEL_TEXT ROM4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>694,-65.5</position>
<gparam>LABEL_TEXT ROM3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>718.5,-55.5</position>
<gparam>LABEL_TEXT ROM5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>718.5,-73.5</position>
<gparam>LABEL_TEXT ROM6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>75</ID>
<type>FF_GND</type>
<position>649.5,-59</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>79</ID>
<type>FF_GND</type>
<position>658,-81.5</position>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>FF_GND</type>
<position>651.5,-81.5</position>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>82</ID>
<type>FF_GND</type>
<position>664.5,-35.5</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>103</ID>
<type>FF_GND</type>
<position>666.5,-35.5</position>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>FF_GND</type>
<position>668.5,-35.5</position>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,692.5</position>
<input>
<ID>IN_0</ID>403 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,687.5</position>
<input>
<ID>IN_0</ID>400 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,682.5</position>
<input>
<ID>IN_0</ID>392 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,677</position>
<input>
<ID>IN_0</ID>391 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,672</position>
<input>
<ID>IN_0</ID>386 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,698</position>
<input>
<ID>IN_0</ID>406 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,667</position>
<input>
<ID>IN_0</ID>225 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_MUX_2x1</type>
<position>1296.5,661.5</position>
<input>
<ID>IN_0</ID>224 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1282.5,671,1282.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_2</name></connection>
<intersection>671 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1282.5,671,1294.5,671</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>1282.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1283.5,676,1283.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_3</name></connection>
<intersection>676 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1283.5,676,1294.5,676</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>1283.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1284.5,681.5,1284.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_4</name></connection>
<intersection>681.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1284.5,681.5,1294.5,681.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>1284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1301.5,685.5,1301.5,698</points>
<intersection>685.5 1</intersection>
<intersection>698 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1301.5,685.5,1316,685.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_7</name></connection>
<intersection>1301.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1298.5,698,1301.5,698</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>1301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1285.5,686.5,1285.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_5</name></connection>
<intersection>686.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1285.5,686.5,1294.5,686.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>1285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1286.5,691.5,1286.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_6</name></connection>
<intersection>691.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1286.5,691.5,1294.5,691.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>1286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1287.5,697,1287.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_7</name></connection>
<intersection>697 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1287.5,697,1294.5,697</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>1287.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1301.5,684.5,1301.5,692.5</points>
<intersection>684.5 2</intersection>
<intersection>692.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1298.5,692.5,1301.5,692.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>1301.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1301.5,684.5,1316,684.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_6</name></connection>
<intersection>1301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>653,-84.5,675,-84.5</points>
<connection>
<GID>20</GID>
<name>SEL_0</name></connection>
<connection>
<GID>24</GID>
<name>SEL_0</name></connection>
<connection>
<GID>25</GID>
<name>SEL_0</name></connection>
<connection>
<GID>26</GID>
<name>SEL_0</name></connection>
<intersection>653 29</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>653,-84.5,653,-62.5</points>
<intersection>-84.5 1</intersection>
<intersection>-62.5 30</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>653,-62.5,696,-62.5</points>
<intersection>653 29</intersection>
<intersection>696 31</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>696,-62.5,696,-61.5</points>
<connection>
<GID>51</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-62.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1280.5,660.5,1280.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>660.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1280.5,660.5,1294.5,660.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>1280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1281.5,666,1281.5,707</points>
<connection>
<GID>195</GID>
<name>OUT_1</name></connection>
<intersection>666 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1281.5,666,1294.5,666</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>1281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>683,-87.5,683,-42.5</points>
<intersection>-87.5 2</intersection>
<intersection>-86 5</intersection>
<intersection>-70 4</intersection>
<intersection>-55 11</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>683,-42.5,689.5,-42.5</points>
<connection>
<GID>50</GID>
<name>ADDRESS_3</name></connection>
<intersection>683 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>650.5,-87.5,683,-87.5</points>
<intersection>650.5 3</intersection>
<intersection>683 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>650.5,-87.5,650.5,-86.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>683,-70,689.5,-70</points>
<connection>
<GID>53</GID>
<name>ADDRESS_3</name></connection>
<intersection>683 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>683,-86,712.5,-86</points>
<intersection>683 0</intersection>
<intersection>690 6</intersection>
<intersection>712.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>690,-88,690,-86</points>
<connection>
<GID>49</GID>
<name>ADDRESS_3</name></connection>
<intersection>-86 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>712.5,-86,712.5,-60.5</points>
<intersection>-86 5</intersection>
<intersection>-78.5 9</intersection>
<intersection>-60.5 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>712.5,-78.5,713.5,-78.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_3</name></connection>
<intersection>712.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>712.5,-60.5,713.5,-60.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_3</name></connection>
<intersection>712.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>683,-55,689.5,-55</points>
<connection>
<GID>51</GID>
<name>ADDRESS_3</name></connection>
<intersection>683 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>684,-91.5,684,-43.5</points>
<intersection>-91.5 5</intersection>
<intersection>-88 2</intersection>
<intersection>-71 4</intersection>
<intersection>-56 13</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>684,-43.5,689.5,-43.5</points>
<connection>
<GID>50</GID>
<name>ADDRESS_2</name></connection>
<intersection>684 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>657,-88,684,-88</points>
<intersection>657 3</intersection>
<intersection>684 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>657,-88,657,-86.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>684,-71,689.5,-71</points>
<connection>
<GID>53</GID>
<name>ADDRESS_2</name></connection>
<intersection>684 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>684,-91.5,688.5,-91.5</points>
<intersection>684 0</intersection>
<intersection>688.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>688.5,-91.5,688.5,-79.5</points>
<intersection>-91.5 5</intersection>
<intersection>-89 10</intersection>
<intersection>-79.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>688.5,-79.5,713.5,-79.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_2</name></connection>
<intersection>688.5 6</intersection>
<intersection>712.5 11</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>688.5,-89,690,-89</points>
<connection>
<GID>49</GID>
<name>ADDRESS_2</name></connection>
<intersection>688.5 6</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>712.5,-79.5,712.5,-61.5</points>
<intersection>-79.5 9</intersection>
<intersection>-61.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>712.5,-61.5,713.5,-61.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_2</name></connection>
<intersection>712.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>684,-56,689.5,-56</points>
<connection>
<GID>51</GID>
<name>ADDRESS_2</name></connection>
<intersection>684 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>684.5,-90.5,684.5,-44.5</points>
<intersection>-90.5 5</intersection>
<intersection>-88.5 2</intersection>
<intersection>-72 4</intersection>
<intersection>-57 11</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>684.5,-44.5,689.5,-44.5</points>
<connection>
<GID>50</GID>
<name>ADDRESS_1</name></connection>
<intersection>684.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>665,-88.5,684.5,-88.5</points>
<intersection>665 3</intersection>
<intersection>684.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>665,-88.5,665,-86.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>684.5,-72,689.5,-72</points>
<connection>
<GID>53</GID>
<name>ADDRESS_1</name></connection>
<intersection>684.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>684.5,-90.5,712.5,-90.5</points>
<intersection>684.5 0</intersection>
<intersection>690 10</intersection>
<intersection>712.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>712.5,-90.5,712.5,-62.5</points>
<intersection>-90.5 5</intersection>
<intersection>-80.5 9</intersection>
<intersection>-62.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>712.5,-62.5,713.5,-62.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_1</name></connection>
<intersection>712.5 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>712.5,-80.5,713.5,-80.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_1</name></connection>
<intersection>712.5 6</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>690,-90.5,690,-90</points>
<connection>
<GID>49</GID>
<name>ADDRESS_1</name></connection>
<intersection>-90.5 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>684.5,-57,689.5,-57</points>
<connection>
<GID>51</GID>
<name>ADDRESS_1</name></connection>
<intersection>684.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>695,-50.5,695,-49</points>
<connection>
<GID>50</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>665,-72.5,665,-50.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>665,-50.5,695,-50.5</points>
<intersection>665 1</intersection>
<intersection>695 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>685.5,-91,685.5,-45.5</points>
<intersection>-91 6</intersection>
<intersection>-89 2</intersection>
<intersection>-73 4</intersection>
<intersection>-58 11</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>685.5,-45.5,689.5,-45.5</points>
<connection>
<GID>50</GID>
<name>ADDRESS_0</name></connection>
<intersection>685.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>672.5,-89,685.5,-89</points>
<intersection>672.5 3</intersection>
<intersection>685.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>672.5,-89,672.5,-86.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>685.5,-73,689.5,-73</points>
<connection>
<GID>53</GID>
<name>ADDRESS_0</name></connection>
<intersection>685.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>685.5,-91,712.5,-91</points>
<connection>
<GID>49</GID>
<name>ADDRESS_0</name></connection>
<intersection>685.5 0</intersection>
<intersection>712.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>712.5,-91,712.5,-63.5</points>
<intersection>-91 6</intersection>
<intersection>-81.5 10</intersection>
<intersection>-63.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>712.5,-63.5,713.5,-63.5</points>
<connection>
<GID>65</GID>
<name>ADDRESS_0</name></connection>
<intersection>712.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>712.5,-81.5,713.5,-81.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_0</name></connection>
<intersection>712.5 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>685.5,-58,689.5,-58</points>
<connection>
<GID>51</GID>
<name>ADDRESS_0</name></connection>
<intersection>685.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>667,-72.5,667,-72.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>55</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666.5,-66.5,666.5,-42.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>-66.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>666,-66.5,666.5,-66.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>666.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>651.5,-80.5,651.5,-79</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>649.5,-80.5,651.5,-80.5</points>
<intersection>649.5 7</intersection>
<intersection>651.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>649.5,-82.5,649.5,-80.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>696,-51.5,696,-49</points>
<connection>
<GID>50</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>671.5,-82.5,671.5,-51.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>671.5,-51.5,696,-51.5</points>
<intersection>671.5 1</intersection>
<intersection>696 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668,-66.5,668,-62</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-62 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>668,-62,695,-62</points>
<intersection>668 0</intersection>
<intersection>695 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>695,-62,695,-61.5</points>
<connection>
<GID>51</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-62 3</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>699.5,-44.5,699.5,-44.5</points>
<connection>
<GID>50</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>699.5,-57,699.5,-57</points>
<connection>
<GID>51</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>699.5,-72,699.5,-72</points>
<connection>
<GID>53</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>700,-90,700,-90</points>
<connection>
<GID>49</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>723.5,-62.5,723.5,-62.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>65</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>723.5,-80.5,723.5,-80.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>650.5,-73,650.5,-66</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<connection>
<GID>68</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654,-73,654,-49</points>
<intersection>-73 4</intersection>
<intersection>-49 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>654,-49,693,-49</points>
<connection>
<GID>50</GID>
<name>DATA_OUT_3</name></connection>
<intersection>654 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>652.5,-73,654,-73</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>654 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>651.5,-60.5,651.5,-60</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>-60.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>693,-61.5,693,-60.5</points>
<connection>
<GID>51</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>651.5,-60.5,693,-60.5</points>
<intersection>651.5 0</intersection>
<intersection>693 1</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>656,-82.5,656,-49.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>694,-49.5,694,-49</points>
<connection>
<GID>50</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>656,-49.5,694,-49.5</points>
<intersection>656 0</intersection>
<intersection>694 1</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664,-82.5,664,-80.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>666,-80.5,666,-78.5</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>664,-80.5,666,-80.5</points>
<intersection>664 0</intersection>
<intersection>666 1</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,-82.5,666,-82.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>673.5,-82.5,673.5,-82.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>649.5,-60,649.5,-60</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>658,-82.5,658,-82.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>651.5,-82.5,651.5,-82.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,-36.5,664.5,-36.5</points>
<connection>
<GID>47</GID>
<name>IN_2</name></connection>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666.5,-36.5,666.5,-36.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-36.5,668.5,-36.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1301.5,683.5,1301.5,687.5</points>
<intersection>683.5 1</intersection>
<intersection>687.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1301.5,683.5,1316,683.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_5</name></connection>
<intersection>1301.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1298.5,687.5,1301.5,687.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>1301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1298.5,682.5,1316,682.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1301.5,677,1301.5,681.5</points>
<intersection>677 2</intersection>
<intersection>681.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1301.5,681.5,1316,681.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_3</name></connection>
<intersection>1301.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1298.5,677,1301.5,677</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>1301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1301.5,672,1301.5,680.5</points>
<intersection>672 1</intersection>
<intersection>680.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1298.5,672,1301.5,672</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>1301.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1301.5,680.5,1316,680.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_2</name></connection>
<intersection>1301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1301.5,667,1301.5,679.5</points>
<intersection>667 1</intersection>
<intersection>679.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1298.5,667,1301.5,667</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>1301.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1301.5,679.5,1316,679.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_1</name></connection>
<intersection>1301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1303,661.5,1303,678.5</points>
<intersection>661.5 2</intersection>
<intersection>678.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1303,678.5,1316,678.5</points>
<connection>
<GID>7</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>7</GID>
<name>DATA_IN_0</name></connection>
<intersection>1303 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1298.5,661.5,1303,661.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>1303 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>96.14,2728.32,1874.14,1810.32</PageViewport>
<gate>
<ID>206</ID>
<type>GA_LED</type>
<position>134.5,49.5</position>
<input>
<ID>N_in3</ID>399 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>GA_LED</type>
<position>137.5,49</position>
<input>
<ID>N_in3</ID>398 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>GA_LED</type>
<position>140.5,49</position>
<input>
<ID>N_in3</ID>397 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>GA_LED</type>
<position>143.5,49</position>
<input>
<ID>N_in3</ID>393 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>EE_VDD</type>
<position>134,58.5</position>
<output>
<ID>OUT_0</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>219</ID>
<type>BB_CLOCK</type>
<position>147,57.5</position>
<output>
<ID>CLK</ID>402 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_REGISTER4</type>
<position>138,56.5</position>
<input>
<ID>IN_0</ID>390 </input>
<input>
<ID>IN_1</ID>389 </input>
<input>
<ID>IN_2</ID>387 </input>
<input>
<ID>IN_3</ID>388 </input>
<output>
<ID>OUT_0</ID>399 </output>
<output>
<ID>OUT_1</ID>398 </output>
<output>
<ID>OUT_2</ID>397 </output>
<output>
<ID>OUT_3</ID>393 </output>
<input>
<ID>clock</ID>401 </input>
<input>
<ID>load</ID>402 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_TOGGLE</type>
<position>137,65.5</position>
<output>
<ID>OUT_0</ID>390 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_TOGGLE</type>
<position>138,63</position>
<output>
<ID>OUT_0</ID>389 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_TOGGLE</type>
<position>139,66</position>
<output>
<ID>OUT_0</ID>387 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_TOGGLE</type>
<position>140,65</position>
<output>
<ID>OUT_0</ID>388 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,60.5,139,64</points>
<connection>
<GID>163</GID>
<name>IN_2</name></connection>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,60.5,140,63</points>
<connection>
<GID>163</GID>
<name>IN_3</name></connection>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,60.5,138,61</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,60.5,137,63.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,51.5,140,52.5</points>
<connection>
<GID>163</GID>
<name>OUT_3</name></connection>
<intersection>51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>143.5,50,143.5,51.5</points>
<connection>
<GID>210</GID>
<name>N_in3</name></connection>
<intersection>51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>140,51.5,143.5,51.5</points>
<intersection>140 0</intersection>
<intersection>143.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,51.5,139,52.5</points>
<connection>
<GID>163</GID>
<name>OUT_2</name></connection>
<intersection>51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>140.5,50,140.5,51.5</points>
<connection>
<GID>208</GID>
<name>N_in3</name></connection>
<intersection>51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>139,51.5,140.5,51.5</points>
<intersection>139 0</intersection>
<intersection>140.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,50,137.5,52.5</points>
<connection>
<GID>207</GID>
<name>N_in3</name></connection>
<intersection>52.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>137.5,52.5,138,52.5</points>
<connection>
<GID>163</GID>
<name>OUT_1</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,50.5,134.5,51.5</points>
<connection>
<GID>206</GID>
<name>N_in3</name></connection>
<intersection>51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>137,51.5,137,52.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134.5,51.5,137,51.5</points>
<intersection>134.5 0</intersection>
<intersection>137 1</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,57.5,134,57.5</points>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<connection>
<GID>163</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,57.5,143,57.5</points>
<connection>
<GID>219</GID>
<name>CLK</name></connection>
<connection>
<GID>163</GID>
<name>load</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-277.392,4102.3,1500.61,3184.3</PageViewport></page 3>
<page 4>
<PageViewport>-277.392,4102.3,1500.61,3184.3</PageViewport></page 4>
<page 5>
<PageViewport>-277.392,4102.3,1500.61,3184.3</PageViewport></page 5>
<page 6>
<PageViewport>-277.392,4102.3,1500.61,3184.3</PageViewport></page 6>
<page 7>
<PageViewport>-277.392,4102.3,1500.61,3184.3</PageViewport></page 7>
<page 8>
<PageViewport>-277.392,4102.3,1500.61,3184.3</PageViewport></page 8>
<page 9>
<PageViewport>-277.392,4102.3,1500.61,3184.3</PageViewport></page 9></circuit>